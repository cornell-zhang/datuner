`timescale 1ps / 1ps
      
module mBnnXcelHLS_v(clk, reset, xcelreq_busy, xcelreq_vld, xcelreq_data, xcelresp_busy, xcelresp_vld, xcelresp_data, memreq_busy, memreq_vld, memreq_data, memresp_busy, memresp_vld, memresp_data);

      input clk;
      input reset;
      input xcelresp_busy;
      input memreq_busy;
      input [159:0] xcelreq_data;
      input [79:0] memresp_data;
      input xcelreq_vld;
      input memresp_vld;
      output xcelreq_busy;
      output memresp_busy;
      output [68:0] xcelresp_data;
      reg [68:0] xcelresp_data;
      output [109:0] memreq_data;
      output xcelresp_vld;
      output memreq_vld;
      reg vld_1;
      reg rdy_1;
      reg vld_0;
      wire rdy_0;
      reg en_0;
      reg en_1;
      reg en_2;
      reg[31:0] bnn_Add_32Ux32U_32U_1_955_in1;
      reg[9:0] bnn_Add_32Ux10U_32U_1_954_in1;
      wire[31:0] bnn_Add_32Ux10U_32U_1_954_out1;
      wire[31:0] bnn_Add_32Ux32U_32U_1_955_out1;
      reg s_reg_870_stage1;
      reg s_reg_870_stage10;
      reg drain3;
      reg cycle1_state2;
      reg[1:0] cycle2_state2;
      wire bnn_And_1Sx1U_1U_4_29_out1;
      wire bnn_And_1Sx1U_1U_4_25_out1;
      reg memreq_m_unacked_req;
      reg xcelresp_m_unacked_req;
      wire bnn_And_1Sx1U_1U_4_8_out1;
      wire bnn_And_1Sx1U_1U_4_4_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_4054_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_4032_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3849_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3827_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3774_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3724_in3;
      wire[1:0] bnn_N_Mux_2_2_3_4_3545_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3541_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3539_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3533_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3532_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3530_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3520_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3519_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3517_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3515_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3505_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3504_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3502_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3501_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3495_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3490_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3489_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3487_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3481_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3476_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3475_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3473_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3467_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3463_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3462_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3460_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3452_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3450_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3449_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_3446_out1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_4_3445_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3444_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3435_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_3434_out1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_4_3433_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3431_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3430_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3428_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3425_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3423_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3416_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3415_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3414_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3412_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3410_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3408_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3407_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3399_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3398_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3396_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3395_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3393_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3383_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3382_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3380_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3368_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3367_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3354_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3351_in3;
      reg[1:0] bnn_N_Mux_2_4_8_4_3341_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3340_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3330_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3328_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_3312_out1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_4_3311_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3303_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3294_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3288_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3285_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3273_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3271_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3257_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3251_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3237_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3223_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3208_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3200_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3186_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3181_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_3171_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3163_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3148_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3132_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3122_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3111_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3101_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3087_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3077_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3061_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3051_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3041_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3034_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3024_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3018_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_3016_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_3009_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3003_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2994_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2992_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2985_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2970_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2968_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2961_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2956_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2945_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2943_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2936_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2929_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2918_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2916_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2912_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2909_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2902_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2891_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2889_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2888_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2882_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2875_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2865_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2864_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2855_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2848_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2840_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2837_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2835_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2828_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2821_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2816_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2810_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2808_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2801_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_2796_out1_slice;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2793_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2782_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2780_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2773_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_2768_out1_slice;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2767_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2766_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2765_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2754_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2752_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2745_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2738_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2727_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2725_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2718_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2711_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2700_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2698_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2694_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2691_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2684_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2673_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2671_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2670_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2664_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2657_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2647_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2646_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2637_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2630_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2622_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2619_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2617_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2610_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2603_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2598_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2592_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2590_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2583_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2576_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2565_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2563_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2556_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2551_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2550_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2549_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2538_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2536_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2529_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2522_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2511_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2509_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2502_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2495_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2484_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2482_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2478_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2475_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2468_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2457_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2455_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2454_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2448_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2441_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2431_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2430_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2421_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2414_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2406_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2403_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2401_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2394_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2386_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2381_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2375_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2373_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2366_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_2361_out1_slice;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2358_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2347_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2345_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2338_out1;
      reg[1:0] bnn_N_Mux_3_2_6_4_2333_out1_slice;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2332_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2331_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2330_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2320_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2319_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2310_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2304_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2297_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2293_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2287_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2281_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2270_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2268_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2267_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_2264_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2261_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2250_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2236_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2225_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2146_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_2145_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_2144_out1;
      wire[1:0] bnn_N_Mux_2_2_3_4_2143_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_2142_out1;
      reg[1:0] bnn_N_Mux_2_4_8_4_2141_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1688_out1_slice;
      reg[1:0] bnn_N_Mux_3_2_6_1_1687_out1_slice;
      reg s_reg_1064_stage1;
      reg s_reg_1045_stage1;
      reg s_reg_1040_stage1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1499_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1499_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1497_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1491_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1490_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1486_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1482_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1478_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1474_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1471_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1469_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1457_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1455_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1423_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1404_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1392_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1368_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1358_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1356_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1346_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1343_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1341_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1334_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1332_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1329_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1327_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1326_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1323_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1321_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1320_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1319_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1318_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1317_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1316_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1314_in2;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1440_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1314_in3;
      reg bnn_N_Mux_2_2_3_4_1308_ctrl1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1308_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1302_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1299_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1296_out1;
      reg bnn_N_Mux_2_2_3_4_1292_ctrl1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1292_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1290_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1287_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1286_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1285_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1284_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1283_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1276_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1275_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1270_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1268_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1265_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1259_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1258_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1256_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1255_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1254_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1253_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1248_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1243_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1242_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1240_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1239_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1231_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1225_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1223_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1222_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1218_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1217_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1205_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1202_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1155_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1140_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1138_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1123_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1122_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1120_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_1107_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1106_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1104_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1103_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1095_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1089_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1087_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1086_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1081_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1078_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1076_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1069_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1066_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1063_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1061_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1060_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1046_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1044_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1043_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1029_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1026_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1015_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_1014_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1000_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_986_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_985_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_974_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_967_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_966_in3;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_963_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_962_out1;
      wire bnn_Not_1U_1U_4_307_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_66_out1;
      wire bnn_NotEQ_7Ux1U_1U_4_65_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_4_960_out1;
      reg s_reg_1069;
      reg s_reg_1065;
      reg s_reg_1062;
      reg s_reg_1055;
      reg s_reg_1051;
      reg s_reg_1049;
      reg s_reg_1045;
      reg s_reg_1042;
      reg s_reg_1040;
      reg s_reg_1038;
      reg s_reg_1037;
      reg[1:0] s_reg_1033;
      reg[31:0] s_reg_1009;
      reg[31:0] s_reg_1010;
      reg[31:0] s_reg_1011;
      reg s_reg_1006;
      reg[31:0] short_addr_conv_out_mi9;
      reg[31:0] short_addr_out_fmap_mi9;
      reg[31:0] short_addr_in_fmap_mi9;
      reg[31:0] short_addr_kh_mi9;
      reg[31:0] s_reg_1003;
      reg[31:0] short_addr_w_mi9;
      reg short_do_max_pool_mi9;
      reg[63:0] short_n_inputs_mi9;
      reg[63:0] s_reg_897;
      reg[1:0] short_width_mode_mi9;
      reg[1:0] s_reg_872;
      /*signed*/reg[1:0] Bline_buffer_97_mi61;
      /*signed*/reg[1:0] Bline_buffer_96_mi61;
      /*signed*/reg[1:0] Bline_buffer_78_mi61;
      /*signed*/reg[1:0] Bline_buffer_77_mi61;
      reg[1:0] s_reg_887;
      reg[31:0] s_reg_1001;
      reg[31:0] s_reg_1008;
      reg[31:0] s_reg_1017;
      reg[31:0] s_reg_1007;
      reg s_reg_907;
      wire bnn_And_1Sx1U_1U_4_33_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_30_out1;
      wire bnn_Not_1U_1U_4_28_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_24_out1;
      wire bnn_And_1Sx1U_1U_4_12_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_9_out1;
      wire bnn_Not_1U_1U_4_7_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_3_out1;
      reg s_reg_1111_stage1;
      reg s_reg_1066_stage1;
      reg s_reg_1063_stage1;
      reg s_reg_1061_stage1;
      reg s_reg_1048_stage1;
      reg s_reg_1044_stage1;
      wire bnn_NotEQ_2Ux1U_1U_4_701_out1;
      wire bnn_OrReduction_5U_1U_4_64_out1;
      wire bnn_Equal_7Ux1U_1U_4_46_out1;
      wire bnn_Equal_7Ux3U_1U_4_45_out1;
      wire bnn_Equal_5Ux4U_1U_4_44_out1;
      wire bnn_Equal_7Ux3U_1U_4_43_out1;
      wire bnn_Equal_7Ux3U_1U_4_42_out1;
      wire bnn_Equal_7Ux3U_1U_4_41_out1;
      wire bnn_Equal_7Ux2U_1U_4_40_out1;
      wire bnn_Equal_7Ux2U_1U_4_39_out1;
      wire[6:0] bnn_Equal_7Ux2U_1U_4_39_in2;
      wire bnn_Equal_5Ux1U_1U_4_38_out1;
      wire[4:0] bnn_Equal_5Ux1U_1U_4_38_in2;
      reg s_reg_1071;
      reg short_popped_go_0_u0_mi9;
      wire bnn_And_1Sx1U_1U_4_67_out1;
      wire bnn_Equal_1Ux1U_1U_1_1_out1;
      wire bnn_Equal_1Ux1U_1U_1_1_1_out1;
      wire[31:0] bnn_N_Mux_32_2_1_4_69_in2;
      wire[63:0] bnn_N_Mux_64_2_2_4_63_in2;
      wire[1:0] bnn_N_Mux_2_2_3_4_62_in2;
      wire bnn_N_Muxb_1_2_18_4_68_in2;
      reg[63:0] bnn_N_MuxB_64_10_5_4_74_out1;
      wire bnn_And_1Sx1U_1U_4_61_out1;
      wire bnn_And_1Sx1U_1U_4_59_out1;
      wire bnn_And_1Sx1U_1U_4_58_out1;
      wire bnn_And_1Sx1U_1U_4_57_out1;
      wire bnn_And_1Sx1U_1U_4_56_out1;
      wire bnn_And_1Sx1U_1U_4_55_out1;
      wire bnn_And_1Sx1U_1U_4_54_out1;
      wire bnn_And_1Sx1U_1U_4_53_out1;
      wire[6:0] bnn_Equal_7Ux1U_1U_4_46_in2;
      reg[31:0] bnn_N_Mux_32_2_1_4_69_out1;
      reg[31:0] bnn_N_Mux_32_2_1_4_70_out1;
      reg[31:0] bnn_N_Mux_32_2_1_4_71_out1;
      reg[31:0] bnn_N_Mux_32_2_1_4_72_out1;
      reg[31:0] bnn_N_Mux_32_2_1_4_73_out1;
      reg[63:0] bnn_N_Mux_64_2_2_4_63_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_62_out1;
      reg bnn_N_Muxb_1_2_18_4_68_out1;
      reg[4:0] global_state_next;
      reg[4:0] global_state;
      reg gs_ctrl599;
      reg[1:0] gs_ctrl74;
      reg[1:0] gs_ctrl23;
      reg gs_ctrl0;
      reg gs_ctrl61;
      reg[1:0] gs_ctrl267;
      reg[1:0] gs_ctrl266;
      reg[1:0] gs_ctrl264;
      reg[1:0] gs_ctrl242;
      reg[1:0] gs_ctrl240;
      reg[1:0] gs_ctrl228;
      reg[1:0] gs_ctrl226;
      reg[1:0] gs_ctrl224;
      reg gs_ctrl222;
      reg gs_ctrl219;
      reg[1:0] gs_ctrl217;
      reg[2:0] gs_ctrl214;
      reg[1:0] gs_ctrl211;
      reg[2:0] gs_ctrl210;
      reg[2:0] gs_ctrl206;
      reg[2:0] gs_ctrl205;
      reg[1:0] gs_ctrl199;
      reg gs_ctrl198;
      reg gs_ctrl105;
      reg[1:0] gs_ctrl196;
      reg[2:0] gs_ctrl820;
      reg gs_ctrl197;
      reg[2:0] gs_ctrl692;
      reg gs_ctrl691;
      reg gs_ctrl690;
      reg gs_ctrl4;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_180_in1_slice;
      wire[2:0] bnn_Add_2Ux2U_3U_4_4427_out1;
      reg[63:0] s_reg_1005;
      wire bnn_GreaterThan_64Ux10U_1U_4_149_out1;
      /*signed*/wire[7:0] bnn_LeftShift_5Sx2U_8S_4_76_out1;
      wire bnn_GreaterThan_32Ux6U_1U_4_179_out1;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r15;
      reg fixed_buffer_0_if_2_wen0_wire;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r15;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r15;
      reg fixed_buffer_0_if_0_wen0_wire;
      reg fixed_buffer_32_if_2_wen0_wire;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r0;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r1;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r2;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r3;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r4;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r5;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r6;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r7;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r8;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r9;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r10;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r11;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r12;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r13;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r14;
      /*signed*/reg[11:0] fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r15;
      reg[3:0] in1_waddr_wire;
      reg[9:0] s_reg_1163;
      reg[9:0] s_reg_1019;
      wire bnn_LessThan_10Ux32U_1U_4_4104_out1;
      reg[6:0] s_reg_1025;
      wire bnn_LessThan_2Ux2U_1U_4_239_out1;
      reg[1:0] bnn_Add_2Ux1U_2U_4_208_in2;
      wire[1:0] bnn_Add_2Ux1U_2U_4_208_out1;
      wire bnn_LessThan_2Ux2U_1U_4_238_out1;
      reg[4:0] s_reg_1032_stage1_slice;
      reg[4:0] s_reg_1029_stage1_slice;
      reg[4:0] s_reg_1031_stage1_slice;
      reg[4:0] s_reg_1021_stage1_slice;
      reg[4:0] s_reg_1030_stage1;
      reg[4:0] s_reg_1027_stage1;
      wire bnn_OrReduction_4U_1U_4_226_out1;
      wire bnn_Equal_4Ux1U_1U_4_225_out1;
      wire bnn_Equal_4Ux2U_1U_4_224_out1;
      wire bnn_Equal_4Ux2U_1U_4_223_out1;
      wire bnn_Equal_4Ux3U_1U_4_222_out1;
      wire bnn_Equal_4Ux3U_1U_4_221_out1;
      wire bnn_Equal_4Ux3U_1U_4_220_out1;
      wire bnn_Equal_4Ux3U_1U_4_219_out1;
      /*signed*/wire[4:0] bnn_Add_5Sx3S_5S_1_211_out1;
      /*signed*/reg[6:0] bnn_Add_7Sx5S_7S_4_195_in2;
      reg[4:0] bnn_Equal_5Ux4U_1U_4_44_in2;
      reg bnn_N_Muxb_1_2_18_4_237_out1;
      reg bnn_N_Muxb_1_2_18_4_236_out1;
      reg bnn_N_Muxb_1_2_18_4_235_out1;
      reg bnn_N_Muxb_1_2_18_4_234_out1;
      reg bnn_N_Muxb_1_2_18_4_233_out1;
      reg bnn_N_Muxb_1_2_18_4_232_out1;
      reg bnn_N_Muxb_1_2_18_4_231_out1;
      reg bnn_N_Muxb_1_2_18_4_229_out1;
      reg bnn_N_Muxb_1_2_18_4_230_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_216_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_215_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_214_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_213_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_212_out1;
      reg[5:0] s_reg_1032;
      reg[5:0] s_reg_1031;
      reg[4:0] s_reg_1030;
      reg[5:0] s_reg_1029;
      reg[3:0] s_reg_1028;
      /*signed*/wire[5:0] bnn_Add_6Sx4S_6S_1_193_out1;
      reg[5:0] s_reg_1021;
      reg[3:0] s_reg_1026;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_180_out1;
      wire[2:0] bnn_N_Mux_3_2_6_4_3446_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_3434_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_3312_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_2796_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_2768_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_2361_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_2333_in2;
      reg[1:0] bnn_N_Mux_2_4_7_4_2177_out1;
      reg[1:0] bnn_N_Mux_2_4_7_4_1921_out1;
      reg[1:0] bnn_N_Mux_2_4_7_4_1919_out1;
      reg[1:0] bnn_N_Mux_2_4_9_4_1834_out1;
      reg[1:0] bnn_N_Mux_2_4_9_4_1832_out1;
      wire[2:0] bnn_N_Mux_3_2_6_4_1640_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_1638_in2;
      wire[2:0] bnn_N_Mux_3_2_6_4_1637_in2;
      reg[1:0] bnn_N_Mux_2_4_7_4_958_out1;
      wire bnn_Not_1U_1U_4_207_out1;
      wire bnn_LessThan_3Ux3U_1U_4_190_out1;
      /*signed*/reg[1:0] Bline_buffer_119_mi61;
      /*signed*/reg[1:0] Bline_buffer_20_mi61;
      reg[2:0] bnn_N_Mux_3_2_6_4_4105_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3019_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2998_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2995_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2974_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2971_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2949_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2946_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2922_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2919_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2895_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2892_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2868_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2865_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2841_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2838_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2814_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2811_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2786_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2783_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2758_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2755_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2731_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2728_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2704_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2701_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2677_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2647_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2623_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2431_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2407_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1328_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1297_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1278_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1079_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1064_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1061_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1044_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1000_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_986_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1482_out1;
      reg[2:0] s_reg_1022;
      /*signed*/reg[7:0] s_reg_1020_stage1_slice;
      reg[9:0] bnn_Add_10Ux1U_10U_4_192_in2;
      wire bnn_LessThan_10Ux32U_1U_4_1576_out1;
      wire[9:0] bnn_Add_10Ux1U_10U_4_192_out1;
      reg s_reg_1112;
      wire bnn_Equal_1Ux1U_1U_1_1_2_out1;
      reg cycle2_state;
      reg drain2;
      reg cycle1_state;
      /*signed*/reg[63:0] bnn_RightShift_64Sx8S_1S_1_228_in2;
      reg[63:0] bnn_N_Mux_64_2_2_1_1636_out1;
      wire bnn_OrReduction_2U_1U_4_241_out1;
      reg s_reg_1078;
      reg[9:0] s_reg_1020;
      reg[9:0] s_reg_1034;
      /*signed*/wire[3:0] bnn_Sub_4Ux1U_4S_4_1538_out1;
      /*signed*/wire[3:0] bnn_Sub_4Ux1U_4S_4_1597_out1;
      reg[9:0] s_reg_1034_stage1;
      /*signed*/wire[11:0] in1_din_wire_31;
      /*signed*/wire[11:0] in1_din_wire_32;
      /*signed*/wire[11:0] in1_din_wire_33;
      /*signed*/wire[11:0] in1_din_wire_34;
      /*signed*/wire[11:0] in1_din_wire_35;
      /*signed*/wire[11:0] in1_din_wire_36;
      /*signed*/wire[11:0] in1_din_wire_37;
      /*signed*/wire[11:0] in1_din_wire_38;
      /*signed*/wire[11:0] in1_din_wire_39;
      /*signed*/wire[11:0] in1_din_wire_40;
      /*signed*/wire[11:0] in1_din_wire_41;
      /*signed*/wire[11:0] in1_din_wire_42;
      /*signed*/wire[11:0] in1_din_wire_43;
      /*signed*/wire[11:0] in1_din_wire_44;
      /*signed*/wire[11:0] in1_din_wire_45;
      /*signed*/wire[11:0] in1_din_wire_46;
      /*signed*/wire[11:0] in1_din_wire_47;
      /*signed*/wire[11:0] in1_din_wire_48;
      reg[3:0] in2_waddr_wire_31;
      reg[3:0] in1_raddr_wire_31;
      /*signed*/wire[11:0] in1_din_wire_49;
      /*signed*/wire[11:0] in1_din_wire_50;
      /*signed*/wire[11:0] in1_din_wire_51;
      /*signed*/wire[11:0] in1_din_wire_52;
      /*signed*/wire[11:0] in1_din_wire_53;
      /*signed*/wire[11:0] in1_din_wire_54;
      /*signed*/wire[11:0] in1_din_wire_55;
      /*signed*/wire[11:0] in1_din_wire_56;
      reg[3:0] in2_waddr_wire_49;
      reg[3:0] in1_raddr_wire_49;
      /*signed*/wire[11:0] in1_din_wire_57;
      reg[3:0] in2_waddr_wire_57;
      reg[3:0] in1_raddr_wire_57;
      /*signed*/wire[11:0] in1_din_wire_58;
      reg[3:0] in2_waddr_wire_58;
      reg[3:0] in1_raddr_wire_58;
      /*signed*/wire[11:0] in1_din_wire_59;
      /*signed*/wire[11:0] in1_din_wire_60;
      /*signed*/wire[11:0] in1_din_wire_61;
      /*signed*/wire[11:0] in1_din_wire_62;
      reg[3:0] in2_waddr_wire_59;
      reg[3:0] in1_raddr_wire_59;
      /*signed*/wire[31:0] bnn_Sub_32Ux1U_32S_1_332_out1;
      wire bnn_LessThanEQ_10Ux33U_1U_4_368_out1;
      reg s_reg_1059_stage1;
      reg[31:0] s_reg_1000;
      /*signed*/wire[11:0] in1_din_wire;
      /*signed*/wire[11:0] in1_din_wire_0;
      /*signed*/wire[11:0] in1_din_wire_1;
      /*signed*/wire[11:0] in1_din_wire_2;
      /*signed*/wire[11:0] in1_din_wire_3;
      /*signed*/wire[11:0] in1_din_wire_4;
      /*signed*/wire[11:0] in1_din_wire_5;
      /*signed*/wire[11:0] in1_din_wire_6;
      /*signed*/wire[11:0] in1_din_wire_7;
      /*signed*/wire[11:0] in1_din_wire_8;
      /*signed*/wire[11:0] in1_din_wire_9;
      /*signed*/wire[11:0] in1_din_wire_10;
      /*signed*/wire[11:0] in1_din_wire_11;
      /*signed*/wire[11:0] in1_din_wire_12;
      /*signed*/wire[11:0] in1_din_wire_13;
      /*signed*/wire[11:0] in1_din_wire_14;
      /*signed*/wire[11:0] in1_din_wire_15;
      /*signed*/wire[11:0] in1_din_wire_16;
      /*signed*/wire[11:0] in1_din_wire_17;
      /*signed*/wire[11:0] in1_din_wire_18;
      /*signed*/wire[11:0] in1_din_wire_19;
      /*signed*/wire[11:0] in1_din_wire_20;
      /*signed*/wire[11:0] in1_din_wire_21;
      /*signed*/wire[11:0] in1_din_wire_22;
      /*signed*/wire[11:0] in1_din_wire_23;
      /*signed*/wire[11:0] in1_din_wire_24;
      /*signed*/wire[11:0] in1_din_wire_25;
      /*signed*/wire[11:0] in1_din_wire_26;
      /*signed*/wire[11:0] in1_din_wire_27;
      /*signed*/wire[11:0] in1_din_wire_28;
      /*signed*/wire[11:0] in1_din_wire_29;
      /*signed*/wire[11:0] in1_din_wire_30;
      wire[3:0] in2_waddr_wire;
      reg[3:0] in1_raddr_wire;
      wire bnn_Equal_2Ux1U_1U_4_78_out1;
      wire bnn_OrReduction_2U_1U_4_77_out1;
      wire bnn_OrReduction_2U_1U_4_3548_out1;
      reg[1:0] bnn_N_Mux_4_2_10_4_80_out1_slice;
      reg[1:0] s_reg_1018_slice;
      wire bnn_OrReduction_2U_1U_4_194_out1;
      wire bnn_OrReduction_2U_1U_4_189_out1;
      wire bnn_OrReduction_2U_1U_4_181_out1;
      reg[3:0] bnn_N_Mux_4_2_11_4_83_out1;
      reg[1:0] s_reg_1004;
      reg[3:0] bnn_N_Mux_4_2_11_4_4100_out1;
      reg[3:0] bnn_N_Mux_4_2_11_4_4099_out1;
      reg[3:0] bnn_N_Mux_4_2_11_4_4098_out1;
      reg[3:0] bnn_N_Mux_4_2_11_4_4090_out1;
      reg[3:0] s_reg_1013;
      /*signed*/reg[2:0] bnn_Add_6Sx4S_6S_1_193_in1_slice;
      /*signed*/reg[5:0] bnn_Add_6Sx4S_6S_1_193_in2;
      wire bnn_LessThan_5Ux32U_1U_4_5204_out1;
      wire bnn_Equal_1Ux1U_1U_1_1_4_out1;
      reg cycle1_state1;
      reg drain;
      reg cycle2_state1;
      /*signed*/reg[11:0] bnn_Mul_30Sx12S_30S_1_191_in1;
      reg[31:0] bnn_Add_32Ux10U_32U_1_954_in2;
      wire bnn_LessThan_5Ux32U_1U_4_5203_out1;
      reg[4:0] s_reg_871_stage1;
      wire bnn_Equal_1Ux1U_1U_1_1_3_out1;
      reg drain1;
      reg cycle2_state0;
      reg cycle1_state0;
      reg cycle3_state;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4988_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4989_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4990_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4991_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4992_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4993_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4994_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4995_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4996_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4997_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4998_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_4999_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5000_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5001_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5002_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5003_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5004_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5005_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5006_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5007_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5008_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5009_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5010_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5011_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5012_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5013_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5014_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5015_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5016_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5017_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5018_in2;
      wire[5:0] bnn_Mod_6Ux32U_7U_4_5019_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4853_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4851_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4848_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4844_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4840_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4836_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4832_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4828_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4824_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4820_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4816_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4812_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4808_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4804_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4800_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4796_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4792_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4788_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4784_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4780_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4776_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4772_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4768_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4764_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4760_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4756_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4752_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4748_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4743_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4737_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4730_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4722_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4713_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4704_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4695_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4686_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4677_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4668_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4659_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4650_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4641_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4632_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4623_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4614_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4605_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4596_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4587_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4578_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4569_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4559_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4549_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4539_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4529_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4519_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4509_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4499_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4489_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4479_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4469_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4459_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4451_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4444_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4438_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4437_in2;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4853_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4851_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4848_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4844_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4840_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4836_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4832_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4828_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4824_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4820_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4816_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4812_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4808_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4804_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4800_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4796_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4792_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4788_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4784_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4780_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4776_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4772_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4768_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4764_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4760_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4756_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4752_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4748_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4743_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4737_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4730_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4722_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4713_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4704_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4695_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4686_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4677_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4668_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4659_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4650_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4641_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4632_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4623_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4614_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4605_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4596_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4587_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4578_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4569_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4559_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4549_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4539_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4529_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4519_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4509_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4499_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4489_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4479_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4469_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4459_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4451_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4444_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4438_out1;
      wire[9:0] bnn_RightShift_10Ux3U_10U_4_4437_out1;
      reg[2:0] s_reg_1012;
      wire bnn_OrReduction_32U_1U_4_4434_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3375_in2;
      reg[5:0] bnn_N_Mux_6_2_12_4_4443_out1;
      wire[6:0] bnn_Mod_2Ux32U_7U_4_4458_out1;
      wire[6:0] bnn_Mod_2Ux32U_7U_4_4450_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4721_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4712_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4703_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4694_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4685_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4676_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4667_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4658_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4649_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4640_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4631_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4622_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4613_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4604_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4595_out1;
      wire[6:0] bnn_Mod_5Ux32U_7U_1_4586_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4577_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4568_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4558_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4548_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4538_out1;
      wire[6:0] bnn_Mod_3Ux32U_7U_4_4468_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4528_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4518_out1;
      wire[6:0] bnn_Mod_3Ux32U_7U_4_4478_out1;
      wire[6:0] bnn_Mod_4Ux32U_7U_4_4508_out1;
      wire[6:0] bnn_Mod_3Ux32U_7U_4_4498_out1;
      wire[6:0] bnn_Mod_3Ux32U_7U_4_4488_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4988_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4989_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4990_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4991_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4992_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4993_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4994_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4995_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4996_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4997_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4998_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_4999_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5000_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5001_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5002_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5003_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5004_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5005_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5006_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5007_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5008_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5009_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5010_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5011_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5012_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5013_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5014_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5015_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5016_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5017_out1;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5018_out1;
      reg[31:0] s_reg_1002;
      wire[6:0] bnn_Mod_6Ux32U_7U_4_5019_out1;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4854_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4852_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4850_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4847_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4843_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4839_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4835_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4831_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4827_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4823_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4819_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4815_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4811_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4807_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4803_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4799_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4795_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4791_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4787_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4783_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4779_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4775_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4771_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4767_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4763_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4759_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4755_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4751_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4747_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4742_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4736_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4729_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4720_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4711_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4702_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4693_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4684_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4675_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4666_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4657_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4648_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4639_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4630_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4621_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4612_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4603_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4594_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4585_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4576_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4567_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4557_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4547_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4537_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4527_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4517_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4507_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4497_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4487_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4477_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4467_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4457_in2;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4449_in2;
      wire[5:0] bnn_LeftShift_1Ux6U_64U_4_4447_in1;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4442_in2;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4441_out1;
      wire[8:0] bnn_LeftShift_9Ux3U_7U_4_4441_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3544_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3544_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3544_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3543_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3543_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3543_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3535_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3535_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3535_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3522_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3522_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3522_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3507_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3507_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3507_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3492_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3492_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3492_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3478_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3478_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3478_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3458_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3458_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3458_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3441_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3441_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3441_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3437_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3437_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3437_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3419_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3419_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3419_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3401_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3401_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3401_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3385_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3385_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3385_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3375_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4442_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3370_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3370_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3370_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3356_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3356_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3356_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3336_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3336_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3336_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3319_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3319_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3319_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3315_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3315_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3315_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3297_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3297_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3297_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3279_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3279_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3279_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3263_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3263_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3263_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3248_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3248_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3248_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3234_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3234_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3234_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3214_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3214_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3214_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3199_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3199_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3199_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3197_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3197_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3197_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3193_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3193_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3193_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3175_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3175_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3175_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3156_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3156_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3156_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3138_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3138_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3138_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3119_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3119_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_3119_in2;
      /*signed*/wire[6:0] bnn_Add_7Sx6U_7S_4_3098_out1;
      reg[5:0] bnn_Add_7Sx6U_7S_4_3098_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4457_out1;
      /*signed*/reg[6:0] bnn_Add_7Sx6U_7S_4_3098_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_4_3070_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_4_3070_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4449_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_4_3070_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2772_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4720_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2772_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2717_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4711_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2717_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2690_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4702_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2690_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2663_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4693_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2663_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2636_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4684_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2636_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2609_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4675_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2609_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2582_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4666_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2582_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2555_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4657_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2555_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2501_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4648_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2501_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2474_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4639_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2474_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2447_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4630_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2447_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2420_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4621_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2420_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2393_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4612_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2393_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2365_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4603_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2365_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2362_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2362_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4594_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2362_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2337_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4585_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2337_in2;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2312_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2312_in1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_2312_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_1526_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4576_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_1526_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_887_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4567_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_887_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_699_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4557_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_699_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_457_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4547_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_457_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_409_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4537_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_409_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_407_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4467_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_407_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_365_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4527_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_365_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_345_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4517_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_345_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_314_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4477_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_314_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_298_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4507_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_298_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_282_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4497_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_282_in2;
      reg[5:0] bnn_Add_6Ux6U_6U_1_274_in1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4487_out1;
      reg[5:0] bnn_Add_6Ux6U_6U_1_274_in2;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4835_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4847_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4729_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4854_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4852_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4763_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4850_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4759_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4843_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4839_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4755_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4771_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4827_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4767_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4823_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4831_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4747_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4815_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_1526_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4751_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4742_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4736_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4811_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4807_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4803_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4799_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4795_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_887_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4791_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4787_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_457_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_409_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4783_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_699_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4819_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4779_out1;
      wire[6:0] bnn_LeftShift_9Ux3U_7U_4_4775_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5148_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5144_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5140_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5136_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5132_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5128_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5124_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5120_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5116_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5112_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5108_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5104_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5100_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5096_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5092_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5088_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5084_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5080_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5076_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5072_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5068_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5064_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5060_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5056_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5052_out1;
      reg[63:0] bnn_N_Mux_64_2_2_4_5048_out1;
      reg[63:0] bnn_N_Mux_64_2_2_4_5044_out1;
      reg[63:0] bnn_N_Mux_64_2_2_4_5040_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5036_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5032_out1;
      reg[63:0] bnn_N_Mux_64_2_2_4_5028_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5024_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4553_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4543_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4533_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4523_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4513_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4503_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4493_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4483_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4473_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4463_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_4746_out1;
      reg[63:0] s_reg_1166;
      reg[63:0] bnn_N_Mux_64_2_2_1_4740_out1;
      reg[63:0] s_reg_1165;
      reg[63:0] bnn_N_Mux_64_2_2_1_4733_out1;
      reg[63:0] s_reg_1164;
      reg[63:0] bnn_N_Mux_64_2_2_1_4725_out1;
      reg[63:0] s_reg_1162;
      reg[63:0] bnn_N_Mux_64_2_2_1_4716_out1;
      reg[63:0] s_reg_1161;
      reg[63:0] bnn_N_Mux_64_2_2_1_4707_out1;
      reg[63:0] s_reg_1160;
      reg[63:0] bnn_N_Mux_64_2_2_1_4698_out1;
      reg[63:0] s_reg_1159;
      reg[63:0] bnn_N_Mux_64_2_2_1_4689_out1;
      reg[63:0] s_reg_1158;
      reg[63:0] bnn_N_Mux_64_2_2_1_4680_out1;
      reg[63:0] s_reg_1157;
      reg[63:0] bnn_N_Mux_64_2_2_1_4671_out1;
      reg[63:0] s_reg_1156;
      reg[63:0] bnn_N_Mux_64_2_2_1_4662_out1;
      reg[63:0] s_reg_1155;
      reg[63:0] bnn_N_Mux_64_2_2_1_4653_out1;
      reg[63:0] s_reg_1154;
      reg[63:0] bnn_N_Mux_64_2_2_1_4644_out1;
      reg[63:0] s_reg_1153;
      reg[63:0] bnn_N_Mux_64_2_2_1_4635_out1;
      reg[63:0] s_reg_1152;
      reg[63:0] bnn_N_Mux_64_2_2_1_4626_out1;
      reg[63:0] s_reg_1151;
      reg[63:0] bnn_N_Mux_64_2_2_1_4617_out1;
      reg[63:0] s_reg_1150;
      reg[63:0] bnn_N_Mux_64_2_2_1_4608_out1;
      reg[63:0] s_reg_1149;
      reg[63:0] bnn_N_Mux_64_2_2_1_4599_out1;
      reg[63:0] s_reg_1148;
      reg[63:0] bnn_N_Mux_64_2_2_1_4590_out1;
      reg[63:0] s_reg_1147;
      reg[63:0] bnn_N_Mux_64_2_2_1_4581_out1;
      reg[63:0] s_reg_1146;
      reg[63:0] bnn_N_Mux_64_2_2_1_4572_out1;
      reg[63:0] s_reg_1145;
      reg[63:0] bnn_N_Mux_64_2_2_1_4563_out1;
      reg[63:0] s_reg_1144;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5200_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5199_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5198_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5197_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5196_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5195_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5194_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5193_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5192_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5191_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5190_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5189_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5188_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5187_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5186_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5185_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5184_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5183_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5182_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5181_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5180_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5179_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5178_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5177_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5176_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5175_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5174_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5173_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5172_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5171_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5170_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5169_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5168_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5167_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5166_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5165_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5164_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5163_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5162_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5161_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5160_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5159_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5158_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5157_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5156_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5155_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5154_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5153_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5152_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5151_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5150_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5149_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5147_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5146_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5143_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5142_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5139_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5138_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5135_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5134_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5131_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5130_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5127_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5126_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5123_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5122_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5119_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5118_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5115_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5114_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5111_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5110_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5107_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5106_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5103_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5102_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5099_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5098_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5095_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5094_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5091_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5090_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5087_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5086_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5083_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5082_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5079_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5078_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5075_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5074_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5071_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5070_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5067_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5066_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5063_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5062_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5059_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_5058_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5055_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_5054_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5051_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_5050_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5047_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5046_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5043_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5042_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5039_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5038_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5035_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5034_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5031_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5030_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5027_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_5026_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_5023_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_5022_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_4_5020_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4741_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4735_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4734_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4727_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4726_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4718_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4717_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4709_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4708_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4700_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4699_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4691_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4690_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4682_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4681_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4673_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4672_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4664_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4663_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4655_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4654_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4646_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4645_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4637_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4636_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4628_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4627_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4619_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4618_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4610_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4609_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4601_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4600_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4592_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4591_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4583_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4582_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4574_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4573_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4565_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4564_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4555_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4554_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4552_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4545_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4544_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4542_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4535_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4534_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4532_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4525_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4524_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4522_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4515_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4514_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4512_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4505_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4504_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4502_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4495_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4494_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4492_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4485_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4484_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4482_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4475_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4474_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4472_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4465_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4464_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_1_4455_out1;
      wire[63:0] bnn_NotBit_64U_64U_4_4454_out1;
      wire[63:0] bnn_LeftShift_1Ux6U_64U_4_4447_out1;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_4562_out1;
      /*signed*/reg[63:0] Boutword_i0_mi87;
      wire bnn_Equal_2Ux2U_1U_4_4460_out1;
      reg[63:0] bnn_N_Mux_64_2_2_1_5202_out1;
      reg[4:0] s_reg_871;
      /*signed*/wire[63:0] bnn_And_64Sx64S_64S_1_5201_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_180_in2;
      /*signed*/wire[6:0] bnn_Add_7Sx5S_7S_4_195_out1;
      reg[5:0] bnn_N_Mux_12_64_13_4_5206_ctrl1;
      reg[31:0] bnn_Add_32Ux32U_32U_1_955_in2;
      reg[11:0] bnn_N_Mux_12_64_13_4_5206_out1;
      /*signed*/reg[11:0] fixed_buffer_0_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_1_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_2_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_3_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_4_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_5_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_6_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_7_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_8_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_9_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_10_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_11_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_12_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_13_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_14_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_15_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_16_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_17_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_18_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_19_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_20_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_21_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_22_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_23_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_24_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_25_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_26_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_27_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_28_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_29_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_30_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_31_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_32_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_33_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_34_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_35_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_36_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_37_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_38_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_39_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_40_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_41_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_42_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_43_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_44_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_45_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_46_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_47_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_48_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_49_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_50_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_51_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_52_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_53_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_54_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_55_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_56_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_57_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_58_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_59_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_60_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_61_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_62_if_1_dout_wire;
      /*signed*/reg[11:0] fixed_buffer_63_if_1_dout_wire;
      reg[1:0] bnn_N_Mux_2_2_3_1_4076_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_4010_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3780_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3730_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3630_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_3407_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3402_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_3393_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3386_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3371_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3357_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2317_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_2293_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2291_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_2270_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2258_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2251_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_2250_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_2244_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2237_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1503_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1490_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1488_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1478_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1476_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1474_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1469_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1461_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1457_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1454_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1452_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1444_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1440_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1437_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1435_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1427_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1423_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1420_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1416_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1413_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1418_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1409_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1407_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1406_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1404_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1402_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1397_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1394_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1392_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1390_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1386_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1379_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1358_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1343_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1327_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1323_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1318_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1316_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1311_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1310_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1306_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1305_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1302_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1301_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1299_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1296_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1295_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1294_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1293_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1290_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1289_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1288_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1287_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1284_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1283_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1258_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1253_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1250_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1242_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1239_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1236_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1229_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1227_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1225_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1222_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1214_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1212_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1210_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1209_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1208_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1207_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1205_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1202_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1196_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1194_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1192_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1191_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1190_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1188_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1186_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1185_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1184_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1176_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1174_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1171_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1170_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1169_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1168_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1165_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1157_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1151_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1148_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1141_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1140_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1134_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1131_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1127_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1126_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1122_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1117_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1114_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1112_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1106_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1103_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1100_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1099_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1098_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1091_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1089_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1086_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1085_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1084_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1074_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1073_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1072_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1071_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1069_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1060_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1058_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1056_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1055_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1054_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1052_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1049_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1048_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1043_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1040_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1038_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1035_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1032_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1031_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1028_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1026_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1020_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1018_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_1014_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1013_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1012_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1011_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1010_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1003_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_1002_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_999_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_998_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_997_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_996_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_993_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_989_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_988_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_985_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_982_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_979_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_977_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_976_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_974_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_971_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_970_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_969_in3;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_968_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_965_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_964_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_963_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_1_962_in1;
      /*signed*/reg[1:0] bnn_Minus_2S_2S_4_960_in1;
      /*signed*/reg[1:0] Bline_buffer_95_mi61;
      /*signed*/reg[1:0] Bline_buffer_94_mi61;
      /*signed*/reg[1:0] Bline_buffer_93_mi61;
      /*signed*/reg[1:0] Bline_buffer_92_mi61;
      /*signed*/reg[1:0] Bline_buffer_91_mi61;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3538_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3537_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3536_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3528_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3527_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3526_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3524_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3523_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3514_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3512_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3511_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3509_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3508_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3499_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3497_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3496_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3494_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3493_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3485_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3483_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3482_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3480_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3479_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3471_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3469_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3468_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3466_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3465_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3456_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3454_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3453_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3443_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3442_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3439_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_3427_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3426_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3424_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3423_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3421_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3420_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3420_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_3411_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3409_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_3409_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_3409_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_3408_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3406_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_3406_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_3406_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3405_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3403_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3402_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3402_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3394_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3392_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3390_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_3390_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_3390_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3389_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3387_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3386_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3386_in2;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3379_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3377_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_3375_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3374_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3373_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3372_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3371_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3371_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3363_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3360_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3359_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3358_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_3358_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_3358_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3357_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3357_in2;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3347_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3346_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3345_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3344_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3343_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3334_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3332_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3331_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3321_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3320_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3317_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3305_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3304_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3302_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3301_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3299_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3298_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3289_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3287_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3286_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3284_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3283_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3281_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3280_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3272_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3270_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3268_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3267_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3265_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3264_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3255_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3253_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3252_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3250_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3249_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3241_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3239_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3238_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3236_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3235_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3227_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3225_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3224_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3222_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3221_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3212_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3210_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3209_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3198_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3195_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3183_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3182_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3180_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3179_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3177_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3176_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3167_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3166_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3165_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3164_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3161_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3160_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3158_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3157_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3150_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3149_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3147_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3145_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3143_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3142_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3140_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3139_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3131_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3130_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3129_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3126_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3124_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3123_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3121_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3120_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_3113_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3112_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3110_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3109_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3108_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3105_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3103_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3102_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3100_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3099_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_3092_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3091_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3089_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3088_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3086_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3085_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3084_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3081_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3079_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3078_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3076_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3075_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_3069_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3068_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_3066_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3065_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3063_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3062_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3060_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3059_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3058_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3055_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_3053_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3052_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_3047_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3046_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_3045_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3044_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_3042_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3041_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_3039_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3038_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3036_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3035_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3033_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3032_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3031_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3028_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3025_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3023_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_3022_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_3020_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_3017_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3016_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_3014_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3013_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3011_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3010_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3008_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3007_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_3006_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_3002_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3001_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3000_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2999_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2996_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2993_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2992_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2990_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2989_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2987_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2986_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2984_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2983_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2982_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2978_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2977_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2975_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2972_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2969_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2968_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2966_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2965_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2963_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2962_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2960_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2959_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2958_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2955_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2954_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2953_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2952_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2950_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2947_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2944_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2943_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2941_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2940_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2938_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2937_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2935_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2934_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2933_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2928_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2927_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2926_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2925_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2923_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2920_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2917_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2916_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2914_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2913_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2911_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2910_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2908_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2907_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2906_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2901_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2900_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2899_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2898_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2896_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2893_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2890_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2889_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2887_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2886_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2884_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2883_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2881_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2880_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2879_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2874_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2873_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2872_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2871_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2869_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2866_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2863_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2862_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2860_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2859_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2857_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2856_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2854_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2853_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2852_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2847_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2846_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2845_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2844_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2842_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2839_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2836_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2835_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2833_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2832_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2830_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2829_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2827_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2826_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2825_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2820_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2819_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2818_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2817_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2815_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2812_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2809_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2808_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2806_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2805_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2803_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2802_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2800_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2799_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2798_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2792_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2791_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2790_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2789_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2787_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2784_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2781_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2780_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2778_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2777_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2775_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2774_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2772_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2771_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2770_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2764_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2763_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2762_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2761_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2759_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2756_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2753_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2752_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2750_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2749_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2747_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2746_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2744_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2743_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2742_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2737_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2736_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2735_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2734_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2732_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2729_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2726_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2725_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2723_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2722_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2720_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2719_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2717_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2716_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2715_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2710_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2709_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2708_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2707_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2705_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2702_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2699_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2698_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2696_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2695_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2693_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2692_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2690_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2689_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2688_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2683_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2682_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2681_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2680_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2678_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2675_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2674_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2672_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2671_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2669_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2668_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2666_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2665_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2663_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2662_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2661_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2656_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2655_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2654_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2653_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2651_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2650_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2648_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2645_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2644_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2642_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2641_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2639_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2638_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2636_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2635_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2634_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2629_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2628_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2627_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2626_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2624_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2621_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2620_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2618_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2617_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2615_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2614_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2612_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2611_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2609_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2608_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2607_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2602_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2601_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2600_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2599_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2597_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2596_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2594_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2593_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2591_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2590_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2588_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2587_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2585_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2584_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2582_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2581_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2580_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2575_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2574_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2573_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2572_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2570_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2569_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2567_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2566_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2564_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2563_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2561_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2560_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2558_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2557_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2555_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2554_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2553_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2548_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2547_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2546_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2545_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2543_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2542_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2540_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2539_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2537_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2536_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2534_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2533_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2531_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2530_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2528_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2527_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2526_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2521_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2520_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2519_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2518_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2516_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2515_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2513_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2512_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2510_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2509_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2507_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2506_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2504_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2503_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2501_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2500_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2499_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2494_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2493_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2492_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2491_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2489_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2488_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2486_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2485_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2483_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2482_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2480_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2479_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2477_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2476_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2474_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2473_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2472_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2467_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2466_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2465_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2464_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2462_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2461_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2459_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2458_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2456_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2455_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2453_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2452_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2450_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2449_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2447_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2446_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2445_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2440_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2439_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2438_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2437_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2435_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2434_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_2432_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2429_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2428_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2426_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2425_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2423_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2422_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2420_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2419_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2418_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2413_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2412_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2411_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2410_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2408_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2405_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2404_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2402_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2401_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2399_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2398_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2396_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2395_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2393_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2392_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2391_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2385_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2384_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2383_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2382_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2380_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2379_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2377_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2376_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2374_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2373_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2371_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2370_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2368_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2367_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2365_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2364_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2363_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2357_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2356_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2355_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2354_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2352_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2351_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2349_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2348_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2346_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2345_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2343_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2342_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2340_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2339_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_2337_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2336_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_2335_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2334_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2329_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2328_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2327_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2326_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2324_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2323_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2321_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2320_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2318_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2317_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2315_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2314_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2311_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2309_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2308_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2303_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2302_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2301_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2300_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2298_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2297_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2295_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2294_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2292_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2291_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_2289_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2288_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2286_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2285_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2280_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2279_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2278_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2277_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2275_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2274_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2272_out1;
      /*signed*/reg[1:0] bnn_Add_4Sx2S_4S_1_2272_in1;
      /*signed*/reg[3:0] bnn_Add_4Sx2S_4S_1_2272_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_2271_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2269_out1;
      /*signed*/reg[1:0] bnn_Add_4Sx2S_4S_1_2269_in1;
      /*signed*/reg[3:0] bnn_Add_4Sx2S_4S_1_2269_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_2268_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2266_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2265_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2260_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2259_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2258_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2257_out1;
      /*signed*/reg[1:0] bnn_Add_2Sx2S_3S_1_2257_in1;
      /*signed*/reg[1:0] bnn_Add_2Sx2S_3S_1_2257_in2;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2255_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2254_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_2252_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2251_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2249_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2248_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2244_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2243_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2242_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2241_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2240_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_2238_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2237_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2235_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2234_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2230_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2229_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2228_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2227_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_2226_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2223_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2220_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2219_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2218_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2216_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_2215_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1635_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1634_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_1542_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1542_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_4032_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1502_in2;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1501_in2;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1500_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_1500_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_3730_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1500_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1499_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1498_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_4_1498_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_4_1498_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1497_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1496_in2;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1495_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1492_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1489_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1489_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1488_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1487_in2;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_4_1485_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1483_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1480_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1479_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1477_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1477_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1476_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1475_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1473_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1470_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1468_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1465_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1464_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1462_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1462_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1461_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1460_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1456_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1454_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1453_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1451_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1448_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1447_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1452_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1445_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1445_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1444_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1443_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1439_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1438_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1436_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1434_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1431_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1430_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1435_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1428_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1428_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1427_out1;
      reg bnn_N_Mux_2_2_3_1_1427_ctrl1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_4_1426_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1422_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1421_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1419_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1417_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1416_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1414_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1413_out1;
      reg bnn_N_Mux_2_2_3_1_1413_ctrl1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1418_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1409_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1408_out1;
      reg bnn_N_Mux_2_2_3_1_1406_ctrl1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1405_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1403_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1400_in2;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1397_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1396_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1395_out1;
      reg bnn_N_Mux_2_2_3_1_1394_ctrl1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1393_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1391_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1391_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1390_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1389_in2;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1386_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1385_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1383_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1382_out1;
      reg bnn_N_Mux_2_2_3_1_1382_ctrl1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1380_out1;
      /*signed*/reg[1:0] bnn_Add_5Sx4S_6S_1_1380_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_3630_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1380_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_1379_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1373_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1366_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1365_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1364_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1363_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1362_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1361_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1360_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1359_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1357_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1356_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1354_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1353_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1352_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1351_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1350_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1349_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1348_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1347_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1345_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1344_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1342_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1341_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1339_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1338_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1337_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1336_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1335_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1334_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_4_1333_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1331_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1330_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1326_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1325_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1324_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1322_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1321_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1315_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_1315_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1314_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_4_1313_in2;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1312_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1311_out1;
      reg bnn_N_Mux_2_2_3_1_1311_ctrl1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1310_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1309_out1;
      /*signed*/reg[1:0] bnn_Add_4Sx2S_5S_4_1309_in1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1486_out1;
      /*signed*/reg[3:0] bnn_Add_4Sx2S_5S_4_1309_in2;
      reg[1:0] bnn_N_Mux_2_2_3_4_1308_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1307_out1;
      reg bnn_N_Mux_2_2_3_1_1306_ctrl1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1305_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1304_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1303_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1300_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1298_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1295_out1;
      reg bnn_N_Mux_2_2_3_1_1294_ctrl1;
      reg bnn_N_Mux_2_2_3_1_1293_ctrl1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_4_1291_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1289_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1288_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1282_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1281_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1279_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1277_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_4_1274_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1273_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1272_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1271_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1270_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1267_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1266_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1265_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1264_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1263_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1262_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1260_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1259_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1257_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1256_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1252_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1251_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1250_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1249_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1247_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1246_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1244_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1243_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1241_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1240_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1238_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1237_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1236_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1235_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1234_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1233_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1232_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1230_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1229_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1227_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1226_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1224_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1223_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1221_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1220_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1219_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1218_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1216_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1215_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1214_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1213_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1212_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1210_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1209_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1208_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1207_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1206_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1204_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1203_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1201_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1200_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1199_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1198_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1197_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1196_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1195_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1194_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1192_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1191_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1190_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1189_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1188_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1187_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1186_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1185_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1184_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1183_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1182_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1181_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1180_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1179_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1178_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1177_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1176_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1175_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1174_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1172_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1171_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1170_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1169_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1168_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1167_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1166_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1165_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1164_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1163_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1162_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1161_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1160_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1159_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1158_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1157_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1156_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1155_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1153_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1152_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1151_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1150_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1149_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1148_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1147_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1146_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1145_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1144_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1143_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1142_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1141_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1139_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1138_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1136_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1135_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1134_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1133_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1132_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1131_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1130_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1129_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1128_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1127_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1126_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1124_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1123_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1121_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1120_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1119_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1118_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1117_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1116_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1115_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1114_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1113_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1112_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1111_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1110_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1108_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1107_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1105_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1104_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1102_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1101_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1100_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1099_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1098_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1097_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1096_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1094_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1093_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1091_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1090_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1088_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1087_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1085_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1084_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1083_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1082_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1080_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1077_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1076_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1074_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1073_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1072_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1071_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1070_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1068_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1067_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1065_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1062_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1059_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1058_out1;
      reg bnn_N_Mux_2_2_3_1_1058_ctrl1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1056_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1055_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1054_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1053_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1052_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1051_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1050_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1049_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1048_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1047_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_1045_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1042_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1041_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1040_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1039_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1038_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1036_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1035_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1033_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1032_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1031_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1030_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1029_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1028_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1027_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1025_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1024_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1023_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1022_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1021_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1020_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1019_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1018_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1017_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1016_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1013_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1012_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1011_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1010_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_1009_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1008_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1007_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1006_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1005_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1004_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1003_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1002_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx3S_4S_1_1001_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_999_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_998_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_997_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_996_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_995_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_994_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_993_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_992_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_991_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_990_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_989_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_988_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_4_987_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_984_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_983_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_982_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_981_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_980_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_979_out1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_978_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_977_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_976_out1;
      reg bnn_N_Mux_2_2_3_1_976_ctrl1;
      /*signed*/wire[2:0] bnn_Add_2Sx2S_3S_1_975_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_973_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_972_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_971_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_970_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_969_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_968_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_967_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_966_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_965_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_964_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1491_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3827_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1471_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1292_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1433_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3780_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1406_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1402_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1467_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1450_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1306_out1;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_216_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_4010_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_216_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_215_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_4_1494_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_215_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_214_in1_slice;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_214_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_213_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_1437_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_213_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx4S_6S_1_212_in1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_4_4060_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx4S_6S_1_212_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx3S_5S_1_211_in1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3516_out1;
      /*signed*/reg[4:0] bnn_Add_5Sx3S_5S_1_211_in2;
      /*signed*/reg[2:0] bnn_Add_5Sx3S_5S_1_209_in1;
      /*signed*/reg[4:0] bnn_Add_5Sx3S_5S_1_209_in2;
      reg[1:0] bnn_N_Mux_2_2_3_1_3349_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_4057_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1301_out1;
      /*signed*/wire[4:0] bnn_Add_5Sx3S_5S_1_209_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1501_out1;
      reg[4:0] s_reg_1143;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1496_out1;
      reg[4:0] s_reg_1142;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1487_out1;
      reg[4:0] s_reg_1141;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1475_out1;
      reg[4:0] s_reg_1140;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1460_out1;
      reg[4:0] s_reg_1139;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1443_out1;
      reg[15:0] s_reg_1138;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1426_out1;
      reg[4:0] s_reg_1137;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1400_out1;
      reg[4:0] s_reg_1136;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1389_out1;
      reg[4:0] s_reg_1135;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1378_out1;
      reg[4:0] s_reg_1134;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1367_out1;
      reg[4:0] s_reg_1133;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1355_out1;
      reg[4:0] s_reg_1132;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1340_out1;
      reg[4:0] s_reg_1131;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1313_out1;
      reg[4:0] s_reg_1130;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1280_out1;
      reg[4:0] s_reg_1129;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1269_out1;
      reg[4:0] s_reg_1128;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1261_out1;
      reg[4:0] s_reg_1127;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1245_out1;
      reg[4:0] s_reg_1126;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1228_out1;
      reg[4:0] s_reg_1125;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1211_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1374_out1;
      reg[4:0] s_reg_1124;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1193_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1371_out1;
      reg[4:0] s_reg_1123;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1173_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_4080_out1;
      reg[4:0] s_reg_1122;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1154_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_4078_out1;
      reg[4:0] s_reg_1121;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1137_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_4076_out1;
      reg[4:0] s_reg_1120;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1125_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1286_out1;
      reg[4:0] s_reg_1119;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1109_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1285_out1;
      reg[4:0] s_reg_1118;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1092_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_4054_out1;
      reg[4:0] s_reg_1117;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1075_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1294_out1;
      reg[4:0] s_reg_1116;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1057_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1384_out1;
      reg[4:0] s_reg_1115;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1037_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3849_out1;
      reg[4:0] s_reg_1114;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_1_1034_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1293_out1;
      reg[4:0] s_reg_1113;
      reg[1:0] bnn_N_Mux_2_2_3_4_1472_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3774_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3724_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1542_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1407_out1;
      /*signed*/wire[1:0] bnn_Minus_2S_2S_1_1503_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1368_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_206_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_1455_out1;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_1_1502_out1;
      /*signed*/wire[3:0] bnn_Add_4Sx2S_4S_1_1372_out1;
      /*signed*/wire[3:0] bnn_Add_3Sx3S_4S_1_1375_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_1369_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1394_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1420_out1;
      reg[4:0] s_reg_1093_stage1_slice;
      reg[4:0] s_reg_1076_stage1_slice;
      reg[4:0] s_reg_1068_stage1_slice;
      /*signed*/reg[6:0] bnn_Add_7Sx4S_7S_1_227_in2;
      /*signed*/reg[4:0] bnn_Add_6Ux6U_6U_1_206_in1_slice;
      reg[5:0] bnn_Add_6Ux6U_6U_1_206_in2;
      /*signed*/reg bnn_LeftShift_2Sx2U_5S_4_75_in2_slice;
      reg[6:0] s_reg_1093;
      reg[6:0] s_reg_1076;
      reg[6:0] s_reg_1068;
      reg s_reg_1088_stage1;
      reg s_reg_1088;
      reg s_reg_1069_stage1;
      wire bnn_N_Mux_3_2_6_4_961_ctrl1;
      wire bnn_N_Mux_3_2_6_4_957_ctrl1;
      reg[1:0] s_reg_998;
      reg[1:0] s_reg_996;
      reg[1:0] s_reg_994;
      reg[1:0] s_reg_992;
      reg[1:0] s_reg_990;
      reg[1:0] s_reg_988;
      reg[1:0] s_reg_986;
      reg[1:0] s_reg_982;
      reg[1:0] s_reg_979;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_961_out1_slice;
      reg[1:0] s_reg_976;
      reg[1:0] s_reg_974;
      reg[1:0] s_reg_971;
      reg[1:0] s_reg_968;
      reg[1:0] s_reg_965;
      reg[1:0] s_reg_962;
      reg[1:0] s_reg_959;
      reg[1:0] s_reg_955;
      reg[1:0] s_reg_949;
      reg[1:0] s_reg_946;
      reg[1:0] s_reg_943;
      reg[1:0] s_reg_941;
      reg[1:0] s_reg_937;
      reg[1:0] s_reg_930;
      reg[1:0] s_reg_927;
      reg[1:0] s_reg_922;
      reg[1:0] s_reg_919;
      reg[1:0] s_reg_914;
      reg[1:0] s_reg_911;
      reg[1:0] s_reg_904;
      reg[1:0] s_reg_900;
      reg[1:0] s_reg_895;
      reg[1:0] s_reg_894;
      reg[1:0] s_reg_890;
      reg[1:0] s_reg_884;
      reg[1:0] s_reg_878;
      reg[1:0] s_reg_873;
      reg s_reg_1094;
      reg s_reg_1087;
      reg s_reg_1077;
      reg[6:0] s_reg_886;
      wire[1:0] bnn_N_Mux_2_2_3_1_2131_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2130_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2130_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2114_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2113_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2113_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2097_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2096_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2096_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2080_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2079_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2079_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2063_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2062_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2062_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2046_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2045_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2045_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2029_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2028_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2028_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2012_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2011_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2011_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2001_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2000_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2000_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1990_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1989_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1989_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1979_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1978_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1978_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1968_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1967_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1967_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1957_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1956_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1956_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1946_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1945_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1945_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1935_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1934_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1934_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1924_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1923_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1923_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1903_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1902_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1902_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1892_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1891_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1891_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1881_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1880_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1880_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1870_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1869_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1869_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1859_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1858_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1858_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1848_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1847_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1847_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1837_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1836_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1836_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1822_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1821_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1821_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1817_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1816_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1816_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1812_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1811_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1811_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1807_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1806_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1806_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1802_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1801_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1801_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1797_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1796_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1796_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1792_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1791_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1791_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1787_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1786_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1786_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_1778_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1777_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1777_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_2198_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_2198_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2197_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_2166_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_2166_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2165_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1914_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1914_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1913_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1529_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1522_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1518_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1518_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1529_out1;
      reg[7:0] s_reg_1096;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1522_out1;
      reg[7:0] s_reg_1089;
      reg[1:0] bnn_N_Mux_3_2_6_1_2180_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_2180_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2179_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2179_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_2154_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_2154_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2153_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2153_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_2148_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_2148_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_2147_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_2147_in1;
      reg[6:0] s_reg_1097;
      reg[4:0] s_reg_1043_stage1;
      reg[4:0] s_reg_1036_stage1;
      reg[4:0] s_reg_1035_stage1;
      reg[4:0] s_reg_1067_stage1_slice;
      reg[4:0] s_reg_1047_stage1;
      reg[4:0] s_reg_1046_stage1_slice;
      reg[5:0] s_reg_1041_stage1_slice;
      reg[4:0] s_reg_1039_stage1;
      reg[5:0] s_reg_1058_stage1_slice;
      /*signed*/reg[4:0] bnn_LeftShift_5Sx2U_8S_4_76_in2;
      reg[6:0] s_reg_1070;
      reg[6:0] s_reg_1067;
      reg[4:0] s_reg_1047;
      reg[6:0] s_reg_1046;
      reg[4:0] s_reg_1043;
      reg[4:0] s_reg_1036;
      reg[4:0] s_reg_1035;
      wire bnn_OrReduction_2U_1U_4_700_out1;
      wire bnn_And_1Sx1U_1U_4_737_out1;
      reg s_reg_1051_stage1;
      reg s_reg_1049_stage1;
      wire bnn_And_1Sx1U_1U_4_1630_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1588_out1;
      wire bnn_Or_1Sx1U_1S_4_1588_in1;
      reg s_reg_1065_stage1;
      wire bnn_And_1Sx1U_1U_4_1587_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1586_out1;
      wire bnn_Or_1Sx1U_1S_4_1586_in1;
      reg s_reg_1062_stage1;
      wire bnn_And_1Sx1U_1U_4_1585_out1;
      reg s_reg_1055_stage1;
      wire bnn_And_1Sx1U_1U_4_1584_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1581_out1;
      wire bnn_Or_1Sx1U_1S_4_1581_in1;
      reg s_reg_1042_stage1;
      wire bnn_And_1Sx1U_1U_4_1580_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1579_out1;
      wire bnn_Or_1Sx1U_1S_4_1579_in1;
      reg s_reg_1038_stage1;
      wire bnn_And_1Sx1U_1U_4_1578_out1;
      reg s_reg_1037_stage1;
      wire bnn_And_1Sx1U_1U_4_1577_out1;
      wire bnn_Or_1Sx1U_1S_4_1519_in1;
      wire bnn_Or_1Sx1U_1S_4_1517_in1;
      wire bnn_Or_1Sx1U_1S_4_1516_in1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1514_out1;
      wire bnn_Or_1Sx1U_1S_4_1514_in1;
      wire bnn_GreaterThan_6Sx4S_1U_4_1513_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1512_out1;
      wire bnn_Or_1Sx1U_1S_4_1512_in1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1511_out1;
      wire bnn_Or_1Sx1U_1S_4_1511_in1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1510_out1;
      wire bnn_Or_1Sx1U_1S_4_1510_in1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1509_out1;
      wire bnn_Or_1Sx1U_1S_4_1509_in1;
      wire bnn_GreaterThan_6Sx4S_1U_4_1508_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1507_out1;
      wire bnn_Or_1Sx1U_1S_4_1507_in1;
      wire bnn_GreaterThan_6Sx4S_1U_4_1506_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1505_out1;
      wire bnn_Or_1Sx1U_1S_4_1505_in1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1504_out1;
      wire bnn_Or_1Sx1U_1S_4_1504_in1;
      wire bnn_And_1Sx1U_1U_4_956_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3545_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3539_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3530_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3517_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3502_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3487_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3473_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3460_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3459_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3447_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3444_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3428_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3412_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3396_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3380_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3365_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3351_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3338_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3337_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3325_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3322_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3306_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3290_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3215_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3274_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_3200_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3258_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3184_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3243_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3168_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3229_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3203_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3151_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3216_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3133_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_959_out1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_3114_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3093_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3071_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1519_out1;
      reg s_reg_1084;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1517_out1;
      reg s_reg_1082;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_1516_out1;
      reg s_reg_1072;
      reg s_reg_1064;
      reg[6:0] s_reg_1058;
      reg[6:0] s_reg_1041;
      reg[4:0] s_reg_1039;
      reg[4:0] s_reg_1027;
      wire bnn_GreaterThan_6Sx4S_1U_4_1515_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_1835_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_99_mi61;
      /*signed*/reg[1:0] Bline_buffer_98_mi61;
      /*signed*/reg[1:0] Bline_buffer_90_mi61;
      /*signed*/reg[1:0] Bline_buffer_69_mi61;
      /*signed*/reg[1:0] Bline_buffer_68_mi61;
      /*signed*/reg[1:0] Bline_buffer_67_mi61;
      /*signed*/reg[1:0] Bline_buffer_66_mi61;
      /*signed*/reg[1:0] Bline_buffer_65_mi61;
      /*signed*/reg[1:0] Bline_buffer_64_mi61;
      /*signed*/reg[1:0] Bline_buffer_63_mi61;
      /*signed*/reg[1:0] Bline_buffer_62_mi61;
      /*signed*/reg[1:0] Bline_buffer_61_mi61;
      /*signed*/reg[1:0] Bline_buffer_60_mi61;
      /*signed*/reg[1:0] Bline_buffer_39_mi61;
      /*signed*/reg[1:0] Bline_buffer_38_mi61;
      /*signed*/reg[1:0] Bline_buffer_37_mi61;
      /*signed*/reg[1:0] Bline_buffer_36_mi61;
      /*signed*/reg[1:0] Bline_buffer_35_mi61;
      /*signed*/reg[1:0] Bline_buffer_34_mi61;
      /*signed*/reg[1:0] Bline_buffer_33_mi61;
      /*signed*/reg[1:0] Bline_buffer_32_mi61;
      /*signed*/reg[1:0] Bline_buffer_31_mi61;
      /*signed*/reg[1:0] Bline_buffer_9_mi61;
      /*signed*/reg[1:0] Bline_buffer_8_mi61;
      /*signed*/reg[1:0] Bline_buffer_7_mi61;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_2178_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_6_mi61;
      /*signed*/reg[1:0] Bline_buffer_5_mi61;
      /*signed*/reg[1:0] Bline_buffer_4_mi61;
      /*signed*/reg[1:0] Bline_buffer_3_mi61;
      /*signed*/reg[1:0] Bline_buffer_2_mi61;
      /*signed*/reg[1:0] Bline_buffer_1_mi61;
      reg s_reg_1044_stage10;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3533_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3520_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3505_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3490_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3476_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3463_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3450_in3;
      reg s_reg_1083_stage1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3415_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3399_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3383_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3368_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3354_in3;
      reg[1:0] bnn_N_Mux_2_2_3_4_3353_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3341_in3;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3328_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3327_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3323_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3313_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3313_in3;
      reg s_reg_1075_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3309_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3308_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3293_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3293_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3292_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3277_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3277_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3276_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3261_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3261_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3260_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3246_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3246_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3245_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3232_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3232_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3231_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3219_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3219_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3218_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3206_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3206_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3205_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3201_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3191_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_3189_out1;
      reg s_reg_1057_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3187_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3172_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3171_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3170_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3154_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3154_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3153_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3136_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3136_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3135_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3117_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3117_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3116_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3096_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3096_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3095_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3074_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3074_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3073_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3050_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3050_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_3049_out1;
      reg s_reg_1056_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_3026_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3026_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2213_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2212_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2211_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2210_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2209_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2207_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2206_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2205_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2204_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2203_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2202_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2201_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2200_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2199_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2195_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2194_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2193_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2192_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2191_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2189_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2188_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2187_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2186_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2185_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2184_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2183_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2182_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2181_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2175_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2174_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2173_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2172_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2171_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2170_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2169_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2168_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2167_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2163_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2162_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2161_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2160_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2159_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2158_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2157_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2156_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2155_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2152_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_2151_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_2150_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2149_out1;
      reg[1:0] bnn_N_Mux_2_2_3_4_2143_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_2141_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2139_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2138_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2137_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2136_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2135_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2135_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2134_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2133_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2132_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2131_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2128_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2127_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2126_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2125_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2124_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2124_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2122_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2121_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2120_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2119_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2118_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2118_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2117_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2116_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2115_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2114_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2111_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2110_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2109_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2108_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2107_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2107_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2105_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2104_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2103_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2102_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2101_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2101_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2100_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2099_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2098_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2097_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2094_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2093_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2092_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2091_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2090_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2090_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2088_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2087_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2086_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2085_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2084_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2084_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2083_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2082_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2081_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2080_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2077_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2076_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2075_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2074_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2073_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2073_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2071_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2070_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2069_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2068_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2067_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2067_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2066_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2065_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2064_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2063_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2060_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2059_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2058_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2057_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2056_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2056_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2054_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2053_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2052_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2051_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2050_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2050_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2049_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2048_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2047_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2046_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2043_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2042_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2041_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2040_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2039_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2039_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2037_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2036_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2035_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2034_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2033_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2033_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2032_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2031_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2030_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2029_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2026_out1;
      reg s_reg_1081_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2025_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2024_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2023_out1;
      reg s_reg_1080_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2022_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2022_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2020_out1;
      reg s_reg_1074_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2019_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2018_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2017_out1;
      reg s_reg_1073_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2016_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2016_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2015_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2014_out1;
      reg s_reg_1079_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2013_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2012_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2009_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2008_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2007_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2006_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2005_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_2005_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_2004_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2003_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_2002_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_2001_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1998_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1997_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1996_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1995_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1994_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1994_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1993_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1992_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1991_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1990_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1987_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1986_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1985_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1984_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1983_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1983_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1982_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1981_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1980_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1979_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1976_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1975_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1974_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1973_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1972_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1972_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1971_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1970_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1969_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1968_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1965_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1964_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1963_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1962_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1961_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1961_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1960_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1959_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1958_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1957_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1954_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1953_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1952_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1951_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1950_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1950_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1949_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1948_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1947_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1946_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1943_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1942_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1941_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1940_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1939_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1939_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1938_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1937_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1936_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1935_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1932_out1;
      reg s_reg_1054_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1931_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1930_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1929_out1;
      reg s_reg_1052_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1928_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1928_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1927_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1926_out1;
      reg s_reg_1085_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1925_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1924_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_1920_out1_slice;
      reg[1:0] bnn_N_Mux_2_2_3_1_1918_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1917_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1916_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1915_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1911_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1910_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1909_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1908_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1907_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1907_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1906_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1905_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1904_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1903_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1900_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1899_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1898_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1897_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1896_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1896_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1895_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1894_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1893_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1892_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1889_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1888_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1887_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1886_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1885_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1885_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1884_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1883_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1882_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1881_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1878_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1877_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1876_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1875_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1874_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1874_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1873_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1872_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1871_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1870_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1867_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1866_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1865_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1864_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1863_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1863_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1862_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1861_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1860_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1859_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1856_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1855_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1854_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1853_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1852_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1852_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1851_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1850_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1849_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1848_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1845_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1844_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1843_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1842_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1841_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1841_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1840_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1839_out1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1838_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1837_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1830_out1;
      reg s_reg_1053_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1829_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1828_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1827_out1;
      reg s_reg_1050_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1826_out1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_1826_in3;
      reg[1:0] bnn_N_Mux_2_2_3_1_1825_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1824_out1;
      reg s_reg_1060_stage1;
      reg[1:0] bnn_N_Mux_2_4_8_1_1823_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1822_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1820_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1819_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1818_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1817_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1815_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1814_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1813_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1812_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1810_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1809_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1808_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1807_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1805_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1804_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1803_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1802_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1800_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1799_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1798_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1797_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1795_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1794_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1793_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1792_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1790_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1789_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1788_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1787_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1785_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_9_4_1784_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1783_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_9_4_1782_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1781_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_1_1780_out1_slice;
      reg[1:0] bnn_N_Mux_2_4_8_1_1779_out1;
      reg[1:0] bnn_N_Mux_2_2_3_1_1778_out1;
      wire bnn_OrReduction_10U_1U_4_1582_out1;
      wire bnn_LessThanEQ_6Sx4S_1U_4_950_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_405_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_394_out1;
      wire bnn_LessThanEQ_5Sx4S_1U_4_358_out1;
      wire bnn_LessThanEQ_6Sx4S_1U_4_348_out1;
      wire bnn_LessThanEQ_5Sx4S_1U_4_338_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_327_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_318_out1;
      wire bnn_LessThanEQ_6Sx4S_1U_4_295_out1;
      wire bnn_LessThanEQ_5Sx4S_1U_4_287_out1;
      wire bnn_LessThanEQ_5Sx4S_1U_4_279_out1;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_957_out1_slice;
      wire bnn_And_1Sx1U_1U_4_315_out1;
      wire bnn_And_1Sx1U_1U_4_952_out1;
      reg s_reg_1111;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_550_out1;
      reg s_reg_1085;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_498_out1;
      reg s_reg_1083;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_487_out1;
      reg s_reg_1081;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_476_out1;
      reg s_reg_1080;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_465_out1;
      reg s_reg_1079;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_453_out1;
      reg s_reg_1075;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_440_out1;
      reg s_reg_1074;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_427_out1;
      reg s_reg_1073;
      /*signed*/wire[4:0] bnn_LeftShift_2Sx2U_5S_4_75_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_454_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_407_out1;
      wire bnn_And_1Sx1U_1U_4_397_out1;
      reg s_reg_1066;
      wire bnn_GreaterThan_6Sx4S_1U_4_503_out1;
      wire bnn_OrReduction_10U_1U_4_280_out1;
      wire bnn_And_1Sx1U_1U_4_386_out1;
      reg s_reg_1063;
      wire bnn_GreaterThan_6Sx4S_1U_4_381_out1;
      wire bnn_And_1Sx1U_1U_4_374_out1;
      reg s_reg_1061;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_370_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_365_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_362_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_360_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_357_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_352_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_350_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_342_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_347_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_340_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_337_out1;
      wire bnn_And_1Sx1U_1U_4_324_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx4S_5S_4_323_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_314_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_308_out1;
      wire bnn_And_1Sx1U_1U_4_305_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx3S_5S_4_304_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_301_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_298_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_294_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx4S_5S_4_290_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_286_out1;
      wire bnn_GreaterThan_6Sx4S_1U_4_278_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx2S_5S_4_276_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx4S_5S_4_272_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_274_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_345_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx3S_5S_4_463_out1;
      /*signed*/wire[4:0] bnn_Add_4Sx4S_5S_4_355_out1;
      wire[5:0] bnn_Add_6Ux6U_6U_1_282_out1;
      reg[1:0] s_reg_977;
      reg[1:0] s_reg_999;
      reg[1:0] s_reg_997;
      reg[1:0] s_reg_984;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_1833_out1_slice;
      reg[1:0] s_reg_995;
      reg[1:0] s_reg_993;
      reg[1:0] s_reg_980;
      reg[1:0] bnn_N_Mux_2_2_3_4_2146_out1;
      reg[1:0] s_reg_991;
      reg[1:0] s_reg_975;
      reg[1:0] bnn_N_Mux_2_2_3_1_2129_out1;
      reg[1:0] s_reg_989;
      reg[1:0] s_reg_972;
      reg[1:0] bnn_N_Mux_2_2_3_1_2112_out1;
      reg[1:0] s_reg_987;
      reg[1:0] s_reg_969;
      reg[1:0] bnn_N_Mux_2_2_3_1_2095_out1;
      reg[1:0] s_reg_985;
      reg[1:0] s_reg_966;
      reg[1:0] bnn_N_Mux_2_2_3_1_2078_out1;
      reg[1:0] s_reg_983;
      reg[1:0] s_reg_981;
      reg[1:0] s_reg_963;
      reg[1:0] bnn_N_Mux_2_2_3_1_2061_out1;
      reg[1:0] s_reg_978;
      reg[1:0] s_reg_960;
      reg[1:0] bnn_N_Mux_2_2_3_1_2044_out1;
      reg[1:0] s_reg_973;
      reg[1:0] s_reg_956;
      reg[1:0] bnn_N_Mux_2_2_3_1_2027_out1;
      reg[1:0] s_reg_950;
      reg[1:0] bnn_N_Mux_2_2_3_1_2214_out1;
      reg[1:0] s_reg_970;
      reg[1:0] s_reg_953;
      reg[1:0] bnn_N_Mux_2_2_3_1_2196_out1;
      reg[1:0] s_reg_967;
      reg[1:0] s_reg_947;
      reg[1:0] bnn_N_Mux_2_2_3_1_2140_out1;
      reg[1:0] s_reg_964;
      reg[1:0] s_reg_942;
      reg[1:0] bnn_N_Mux_2_2_3_1_2123_out1;
      reg[1:0] s_reg_961;
      reg[1:0] s_reg_938;
      reg[1:0] bnn_N_Mux_2_2_3_1_2106_out1;
      reg[1:0] s_reg_958;
      reg[1:0] s_reg_931;
      reg[1:0] bnn_N_Mux_2_2_3_1_2089_out1;
      reg[1:0] s_reg_954;
      reg[1:0] s_reg_923;
      reg[1:0] bnn_N_Mux_2_2_3_1_2072_out1;
      reg[1:0] s_reg_952;
      reg[1:0] s_reg_948;
      reg[1:0] s_reg_915;
      reg[1:0] bnn_N_Mux_2_2_3_1_2055_out1;
      reg[1:0] s_reg_945;
      reg[1:0] s_reg_906;
      reg[1:0] bnn_N_Mux_2_2_3_1_2038_out1;
      reg[1:0] s_reg_940;
      reg[1:0] s_reg_896;
      reg[1:0] bnn_N_Mux_2_2_3_1_2021_out1;
      reg[1:0] s_reg_905;
      reg[1:0] bnn_N_Mux_2_2_3_1_2208_out1;
      reg[1:0] s_reg_936;
      reg[1:0] s_reg_935;
      reg[1:0] bnn_N_Mux_2_2_3_1_2190_out1;
      reg[1:0] s_reg_929;
      reg[1:0] s_reg_928;
      reg[1:0] bnn_N_Mux_2_2_3_1_2010_out1;
      reg[1:0] s_reg_921;
      reg[1:0] s_reg_920;
      reg[1:0] bnn_N_Mux_2_2_3_1_1999_out1;
      reg[1:0] s_reg_913;
      reg[1:0] s_reg_912;
      reg[1:0] bnn_N_Mux_2_2_3_1_1988_out1;
      reg[1:0] s_reg_903;
      reg[1:0] s_reg_901;
      reg[1:0] bnn_N_Mux_2_2_3_1_1977_out1;
      reg[1:0] s_reg_893;
      reg[1:0] s_reg_892;
      reg[1:0] bnn_N_Mux_2_2_3_1_1966_out1;
      reg[1:0] s_reg_934;
      reg[1:0] s_reg_902;
      reg[1:0] s_reg_885;
      reg[1:0] bnn_N_Mux_2_2_3_1_1955_out1;
      reg[1:0] s_reg_926;
      reg[1:0] s_reg_880;
      reg[1:0] bnn_N_Mux_2_2_3_1_1944_out1;
      reg[1:0] s_reg_918;
      reg[1:0] s_reg_879;
      reg[1:0] bnn_N_Mux_2_2_3_1_1933_out1;
      /*signed*/reg[1:0] Bline_buffer_30_mi61;
      reg[1:0] s_reg_891;
      reg[1:0] bnn_N_Mux_2_2_3_1_2176_out1;
      reg[1:0] s_reg_910;
      reg[1:0] s_reg_933;
      reg[1:0] bnn_N_Mux_2_2_3_1_2164_out1;
      reg[1:0] s_reg_899;
      reg[1:0] s_reg_925;
      reg[1:0] bnn_N_Mux_2_2_3_1_1912_out1;
      reg[1:0] s_reg_889;
      reg[1:0] s_reg_917;
      reg[1:0] bnn_N_Mux_2_2_3_1_1901_out1;
      reg[1:0] s_reg_883;
      reg[1:0] s_reg_882;
      reg[1:0] s_reg_909;
      reg[1:0] bnn_N_Mux_2_2_3_1_1890_out1;
      reg[1:0] s_reg_877;
      reg[1:0] s_reg_898;
      reg[1:0] bnn_N_Mux_2_2_3_1_1879_out1;
      reg[1:0] s_reg_876;
      reg[1:0] s_reg_888;
      reg[1:0] bnn_N_Mux_2_2_3_1_1868_out1;
      reg[1:0] s_reg_881;
      reg[1:0] bnn_N_Mux_2_2_3_1_1857_out1;
      reg[1:0] s_reg_875;
      reg[1:0] bnn_N_Mux_2_2_3_1_1846_out1;
      reg[6:0] s_reg_874;
      reg[1:0] bnn_N_Mux_2_2_3_1_1831_out1;
      /*signed*/reg[1:0] Bline_buffer_0_mi61;
      /*signed*/reg[1:0] bnn_N_Mux_3_2_6_4_1922_out1_slice;
      reg s_reg_1044_stage2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3540_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3540_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3531_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3531_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3518_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3518_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3503_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3503_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3488_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3488_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3474_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3474_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3461_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3461_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3448_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3448_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3429_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3429_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3413_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3413_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3397_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3397_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3381_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3381_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3366_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3366_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3365_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3339_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3339_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3338_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3326_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3326_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3322_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3307_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3307_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3306_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3291_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3291_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3290_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3275_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3275_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3274_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3259_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3259_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3258_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3244_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3244_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3243_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3230_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3230_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3229_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3217_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3217_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3216_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3204_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3204_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3185_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3185_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3184_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3169_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3169_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3168_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3152_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3152_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3151_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3134_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3134_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3133_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3115_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3115_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3114_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3094_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3094_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3093_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3072_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3072_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_3071_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3048_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3048_in1;
      wire[1:0] bnn_N_Mux_2_2_3_1_2140_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2137_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2134_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2129_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2126_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2123_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2120_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2117_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2112_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2109_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2106_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2103_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2100_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2095_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2092_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2089_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2086_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2083_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2078_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2075_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2072_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2069_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2066_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2061_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2058_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2055_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2052_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2049_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2044_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2041_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2038_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2035_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2032_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2027_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2024_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2021_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2018_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2015_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2010_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2007_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_2004_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1999_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1996_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1993_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1988_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1985_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1982_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1977_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1974_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1971_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1966_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1963_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1960_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1955_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1952_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1949_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1944_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1941_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1938_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1933_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1930_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1927_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1912_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1909_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1906_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1901_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1898_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1895_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1890_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1887_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1884_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1879_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1876_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1873_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1868_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1865_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1862_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1857_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1854_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1851_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1846_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1843_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1840_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1831_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1828_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1825_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1820_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1815_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1810_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1805_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1800_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1795_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1790_in3;
      wire[1:0] bnn_N_Mux_2_2_3_1_1781_in3;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_1754_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_1754_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1753_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1753_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1752_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1752_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1751_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1751_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1750_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1750_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1749_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1749_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1748_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1748_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1747_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1747_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1746_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1746_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1745_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1745_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1744_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1744_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1743_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1743_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1742_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1742_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1741_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1741_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1740_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1740_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1739_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1739_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1738_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1738_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1737_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1737_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1736_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1736_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1735_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1735_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1734_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1734_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1733_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1733_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1732_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1732_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1731_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1731_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_1730_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_1730_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1729_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1729_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1728_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1728_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1727_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1727_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1726_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1726_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1725_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1725_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1724_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1724_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1723_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1723_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1722_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1722_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1721_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1721_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1720_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1720_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1719_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1719_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1718_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1718_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1717_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1717_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1716_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1716_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1715_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1715_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1714_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1714_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1713_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1713_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1712_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1712_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1711_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1711_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1710_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1710_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1709_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1709_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1708_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1708_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1707_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1707_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1706_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1706_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1705_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1705_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1704_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1704_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1703_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1703_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1702_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1702_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1701_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1701_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1700_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1700_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1699_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1699_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1696_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1696_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1695_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1695_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1694_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1694_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1693_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1693_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1692_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1692_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1691_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1691_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1690_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1690_in1;
      /*signed*/wire bnn_RightShift_64Sx7S_1S_1_1689_out1;
      /*signed*/wire[6:0] bnn_RightShift_64Sx7S_1S_1_1689_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_1674_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_1674_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1673_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1673_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1672_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1672_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1671_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1671_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1670_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1670_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1669_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1669_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1668_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1668_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1667_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1667_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1666_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1666_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1665_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1665_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1664_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1664_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1663_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1663_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1662_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1662_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1661_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1661_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1660_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1660_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1659_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1659_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1658_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1658_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1657_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1657_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1656_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1656_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1655_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1655_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1654_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1654_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1653_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1653_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1652_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1652_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1651_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1651_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_1650_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_1650_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1649_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1649_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1648_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1648_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1647_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1647_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1646_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1646_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1645_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1645_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1644_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1644_in1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1643_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1643_in1;
      /*signed*/reg[7:0] bnn_RightShift_64Sx8S_1S_1_228_in1;
      /*signed*/reg[1:0] Bline_buffer_108_mi61;
      /*signed*/reg[1:0] Bline_buffer_107_mi61;
      /*signed*/reg[1:0] Bline_buffer_106_mi61;
      /*signed*/reg[1:0] Bline_buffer_105_mi61;
      /*signed*/reg[1:0] Bline_buffer_104_mi61;
      /*signed*/reg[1:0] Bline_buffer_103_mi61;
      /*signed*/reg[1:0] Bline_buffer_102_mi61;
      /*signed*/reg[1:0] Bline_buffer_101_mi61;
      /*signed*/reg[1:0] Bline_buffer_76_mi61;
      /*signed*/reg[1:0] Bline_buffer_75_mi61;
      /*signed*/reg[1:0] Bline_buffer_74_mi61;
      /*signed*/reg[1:0] Bline_buffer_73_mi61;
      /*signed*/reg[1:0] Bline_buffer_72_mi61;
      /*signed*/reg[1:0] Bline_buffer_71_mi61;
      /*signed*/reg[1:0] Bline_buffer_48_mi61;
      /*signed*/reg[1:0] Bline_buffer_47_mi61;
      /*signed*/reg[1:0] Bline_buffer_46_mi61;
      /*signed*/reg[1:0] Bline_buffer_45_mi61;
      /*signed*/reg[1:0] Bline_buffer_44_mi61;
      /*signed*/reg[1:0] Bline_buffer_43_mi61;
      /*signed*/reg[1:0] Bline_buffer_42_mi61;
      /*signed*/reg[1:0] Bline_buffer_41_mi61;
      /*signed*/reg[1:0] Bline_buffer_18_mi61;
      /*signed*/reg[1:0] Bline_buffer_17_mi61;
      /*signed*/reg[1:0] Bline_buffer_16_mi61;
      /*signed*/reg[1:0] Bline_buffer_15_mi61;
      /*signed*/reg[1:0] Bline_buffer_14_mi61;
      /*signed*/reg[1:0] Bline_buffer_13_mi61;
      /*signed*/reg[1:0] Bline_buffer_12_mi61;
      /*signed*/reg[1:0] Bline_buffer_11_mi61;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3417_out1;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3295_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_3190_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_3190_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3173_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1776_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1776_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1775_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1772_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1772_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1771_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1768_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1768_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1767_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1764_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1764_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1763_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1760_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1760_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1759_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1698_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1698_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1697_out1;
      wire[2:0] bnn_N_Mux_3_2_6_1_1688_in2;
      reg[1:0] bnn_N_Mux_3_2_6_1_1686_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1686_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1685_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1682_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1682_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1681_out1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1678_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1678_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1677_out1;
      wire[2:0] bnn_N_Mux_3_2_6_1_1642_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1619_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1619_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1610_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1610_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1606_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1606_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1600_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1600_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1596_out1;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1596_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1540_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1536_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1533_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1531_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1527_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1525_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1520_in2;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1540_out1;
      reg[7:0] s_reg_1105;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1536_out1;
      reg[7:0] s_reg_1103;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1533_out1;
      reg[7:0] s_reg_1100;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1531_out1;
      reg[7:0] s_reg_1098;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1527_out1;
      reg[7:0] s_reg_1092;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1525_out1;
      reg[7:0] s_reg_1090;
      /*signed*/wire[7:0] bnn_Sub_8Sx2S_8S_4_1520_out1;
      reg[7:0] s_reg_1086;
      reg[1:0] bnn_N_Mux_3_2_6_1_1642_out1_slice;
      reg[1:0] bnn_N_Mux_3_2_6_4_1638_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_100_mi61;
      /*signed*/reg[1:0] Bline_buffer_70_mi61;
      reg[1:0] bnn_N_Mux_3_2_6_4_1640_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_40_mi61;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_4_3432_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_4_3432_in1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_4_3431_in3;
      reg[1:0] bnn_N_Mux_3_2_6_1_3324_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_3324_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3310_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3310_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_3202_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_3202_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_3188_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_3188_in1;
      /*signed*/wire[1:0] bnn_N_Mux_2_4_8_1_3187_in3;
      reg[1:0] bnn_N_Mux_3_2_6_1_1774_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1774_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1773_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1773_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1770_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1770_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1769_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1769_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1766_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1766_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1765_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1765_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1762_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1762_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1761_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1761_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1758_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1758_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1757_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1757_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1756_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1756_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1755_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1755_in1;
      wire[2:0] bnn_N_Mux_3_2_6_1_1687_in2;
      reg[1:0] bnn_N_Mux_3_2_6_1_1684_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1684_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1683_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1683_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1680_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1680_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1679_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1679_in1;
      reg[1:0] bnn_N_Mux_3_2_6_1_1676_out1_slice;
      wire[2:0] bnn_N_Mux_3_2_6_1_1676_in2;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_1675_out1;
      /*signed*/wire[7:0] bnn_RightShift_64Sx8S_1S_1_1675_in1;
      wire[2:0] bnn_N_Mux_3_2_6_1_1641_in2;
      wire[2:0] bnn_N_Mux_3_2_6_1_1639_in2;
      /*signed*/reg[1:0] bnn_Add_7Sx4S_7S_1_227_in1_slice;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1565_out1;
      reg[4:0] s_reg_1110;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1556_out1;
      reg[4:0] s_reg_1109;
      /*signed*/wire[5:0] bnn_Add_5Sx4S_6S_4_1552_out1;
      reg[4:0] s_reg_1108;
      /*signed*/wire[6:0] bnn_Add_7Sx4S_7S_1_227_out1;
      reg[6:0] s_reg_1107;
      reg[6:0] s_reg_1106;
      reg[6:0] s_reg_1104;
      reg[6:0] s_reg_1102;
      reg[6:0] s_reg_1101;
      reg[4:0] s_reg_1099;
      reg[6:0] s_reg_1095;
      reg[6:0] s_reg_1091;
      reg[1:0] bnn_N_Mux_3_2_6_1_1641_out1_slice;
      reg[1:0] bnn_N_Mux_3_2_6_4_1637_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_79_mi61;
      /*signed*/reg[1:0] Bline_buffer_49_mi61;
      reg[1:0] bnn_N_Mux_3_2_6_1_1639_out1_slice;
      /*signed*/reg[1:0] Bline_buffer_19_mi61;
      reg memreq_m_req_m_trig_req;
      reg xcelresp_m_req_m_trig_req;
      reg memreq_m_req_m_prev_trig_req;
      reg xcelresp_m_req_m_prev_trig_req;
      wire bnn_Not_1U_1U_4_23_out1;
      wire bnn_Not_1U_1U_4_19_out1;
      reg iostall_1;
      reg[159:0] bnn_N_MuxB_160_2_0_4_37_out1;
      reg memresp_m_busy_req_0;
      reg xcelreq_m_busy_req_0;
      wire bnn_Not_1U_1U_4_10_out1;
      wire bnn_Not_1U_1U_4_31_out1;
      reg memresp_m_stall_reg_full;
      reg xcelreq_m_stall_reg_full;
      reg xcelreq_m_stalling;
      reg stall0;
      reg[63:0] memresp_m_stall_reg_slice;
      reg[159:0] xcelreq_m_stall_reg;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_27_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_6_out1;
      reg bnn_N_Muxb_1_2_18_4_2_out1;
      reg memresp_m_unvalidated_req;
      reg bnn_N_Muxb_1_2_18_4_1_out1;
      reg xcelreq_m_unvalidated_req;
      /*signed*/wire bnn_RightShift_64Sx8S_1S_1_228_out1;
      reg s_reg_957;
      reg s_reg_951;
      reg s_reg_944;
      reg s_reg_939;
      reg s_reg_932;
      reg s_reg_924;
      reg s_reg_916;
      reg s_reg_908;
      wire bnn_Not_1U_1U_4_32_out1;
      wire bnn_And_1Sx1U_1U_4_34_out1;
      wire bnn_Not_1U_1U_4_11_out1;
      wire bnn_And_1Sx1U_1U_4_13_out1;
      wire bnn_And_1Sx1U_1U_4_35_out1;
      wire bnn_And_1Sx1U_1U_4_14_out1;
      wire bnn_N_Mux_64_2_2_1_4746_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4740_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4733_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4725_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4716_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4707_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4698_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4689_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4680_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4671_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4662_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4653_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4644_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4635_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4626_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4617_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4608_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4599_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4590_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4581_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4572_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4563_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4553_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4543_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4533_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4523_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4513_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4503_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4493_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4483_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4473_ctrl1;
      wire bnn_N_Mux_64_2_2_1_4463_ctrl1;
      reg s_reg_1060;
      reg s_reg_1059;
      reg s_reg_1057;
      reg s_reg_1056;
      reg s_reg_1054;
      reg s_reg_1053;
      reg s_reg_1052;
      reg s_reg_1050;
      reg s_reg_1048;
      reg s_reg_1044;
      reg s_reg_1024;
      reg s_reg_1023;
      reg s_reg_1016;
      reg s_reg_1015;
      reg s_reg_1014;
      reg s_reg_870;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3547_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3546_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3542_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3534_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3521_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3506_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3491_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3477_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3464_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3451_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3436_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3418_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3400_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3384_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3369_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3355_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3342_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3329_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3314_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3296_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3278_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3262_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3247_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3233_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3220_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3207_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3192_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3174_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3162_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3155_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3146_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3137_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3128_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3118_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3107_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3097_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3083_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3057_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3030_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_3005_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2981_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2957_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2932_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2905_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2878_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2851_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2824_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2797_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2769_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2741_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2714_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2687_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2660_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2633_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2606_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2579_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2552_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2525_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2498_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2471_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2444_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2417_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2390_in2;
      /*signed*/reg[16:0] bnn_Add_17Sx16S_17S_1_2389_in2;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3547_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3546_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3542_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3534_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3521_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3506_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3491_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3477_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3464_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3451_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3436_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3418_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3400_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3384_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3369_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3355_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3342_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3329_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3314_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3296_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3278_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3262_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3247_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3233_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3220_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3207_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3192_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3174_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3162_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3155_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3146_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3137_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3128_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3118_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3107_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3097_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3083_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3057_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3030_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_3005_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2981_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2957_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2932_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2905_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2878_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2851_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2824_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2797_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2769_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2741_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2714_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2687_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2660_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2633_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2606_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2579_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2552_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2525_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2498_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2471_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2444_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2417_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2390_in1;
      /*signed*/reg[15:0] bnn_Add_17Sx16S_17S_1_2389_in1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3146_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3128_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3107_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3083_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3057_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3030_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3005_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2981_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2957_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2932_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2905_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2878_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2851_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2824_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2797_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2769_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2741_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2714_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2687_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2660_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2633_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2606_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2579_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2552_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2525_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2498_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2471_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2444_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2417_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2390_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3547_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3546_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3542_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3534_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3521_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3506_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3491_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3477_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3464_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3451_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3436_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3418_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3400_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3384_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3369_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3355_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3342_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3329_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3233_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3220_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3207_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3192_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3174_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3155_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3137_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3097_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3296_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3262_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3247_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3278_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3314_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3118_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_3162_out1;
      /*signed*/wire[16:0] bnn_Add_17Sx16S_17S_1_2389_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4706_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4697_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4688_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4679_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4670_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4661_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4652_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4643_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4634_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4625_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4616_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4607_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4598_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4589_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4580_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4571_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4561_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4551_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4436_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4462_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4440_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4453_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4446_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4541_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4531_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4521_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4511_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4501_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4430_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4491_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4846_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4481_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4842_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4433_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4838_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4471_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4834_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4830_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4826_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4822_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4818_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4814_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4810_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4806_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4802_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4798_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4794_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4790_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4786_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4782_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4778_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4774_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4770_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4766_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4762_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4758_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4754_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4750_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4745_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4739_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4732_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4724_out1;
      /*signed*/wire[18:0] bnn_Mul_16Sx12S_19S_4_4715_out1;
      /*signed*/reg[29:0] bnn_Mul_30Sx12S_30S_1_191_in2;
      /*signed*/wire[29:0] bnn_Mul_30Sx12S_30S_1_191_out1;
      reg iostall_2;
      reg[96:0] memreq_data_slice;
      wire bnn_Xor_1Ux1U_1U_4_20_out1;
      wire bnn_Xor_1Ux1U_1U_4_16_out1;
      wire bnn_And_1Sx1U_1U_4_18_out1;
      wire bnn_And_1Sx1U_1U_4_22_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_21_out1;
      /*signed*/wire bnn_Or_1Sx1U_1S_4_17_out1;

         // resource: bnn_fixed_buffer_63_regbank
         always @(in1_raddr_wire_59 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r0 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r1 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r2 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r3 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r4 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r5 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r6 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r7 or 
fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r8
          or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r9 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r10 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r11 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r12 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r13 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r14 or fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r15)
          begin :fixed_buffer_63_inst
            case (in1_raddr_wire_59) 

               4'd00: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_63_if_1_dout_wire = fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_63_regbank  instance: fixed_buffer_63_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd15) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r15 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd14) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r14 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd13) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r13 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd12) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r12 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd11) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r11 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd10) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r10 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd09) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r9 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd08) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r8 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd07) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r7 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd06) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r6 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd05) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r5 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd04) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r4 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd03) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r3 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd02) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r2 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd01) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r1 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_63_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_59)) begin
                  fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r0 <= in1_din_wire_62;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_63_inst_bnn_fixed_buffer_63_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_62_regbank
         always @(in1_raddr_wire_59 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r0 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r1 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r2 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r3 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r4 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r5 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r6 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r7 or 
fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r8
          or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r9 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r10 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r11 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r12 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r13 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r14 or fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r15)
          begin :fixed_buffer_62_inst
            case (in1_raddr_wire_59) 

               4'd00: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_62_if_1_dout_wire = fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_62_regbank  instance: fixed_buffer_62_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd15) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r15 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd14) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r14 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd13) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r13 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd12) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r12 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd11) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r11 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd10) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r10 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd09) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r9 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd08) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r8 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd07) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r7 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd06) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r6 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd05) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r5 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd04) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r4 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd03) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r3 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd02) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r2 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd01) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r1 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_62_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_59)) begin
                  fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r0 <= in1_din_wire_61;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_62_inst_bnn_fixed_buffer_62_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_61_regbank
         always @(in1_raddr_wire_59 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r0 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r1 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r2 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r3 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r4 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r5 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r6 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r7 or 
fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r8
          or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r9 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r10 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r11 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r12 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r13 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r14 or fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r15)
          begin :fixed_buffer_61_inst
            case (in1_raddr_wire_59) 

               4'd00: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_61_if_1_dout_wire = fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_61_regbank  instance: fixed_buffer_61_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd15) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r15 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd14) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r14 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd13) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r13 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd12) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r12 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd11) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r11 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd10) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r10 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd09) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r9 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd08) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r8 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd07) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r7 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd06) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r6 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd05) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r5 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd04) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r4 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd03) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r3 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd02) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r2 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd01) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r1 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_61_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_59)) begin
                  fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r0 <= in1_din_wire_60;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_61_inst_bnn_fixed_buffer_61_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_60_regbank
         always @(in1_raddr_wire_59 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r0 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r1 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r2 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r3 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r4 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r5 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r6 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r7 or 
fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r8
          or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r9 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r10 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r11 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r12 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r13 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r14 or fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r15)
          begin :fixed_buffer_60_inst
            case (in1_raddr_wire_59) 

               4'd00: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_60_if_1_dout_wire = fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_60_regbank  instance: fixed_buffer_60_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd15) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r15 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd14) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r14 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd13) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r13 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd12) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r12 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd11) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r11 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd10) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r10 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd09) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r9 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd08) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r8 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd07) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r7 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd06) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r6 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd05) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r5 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd04) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r4 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd03) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r3 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd02) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r2 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_59 == 4'd01) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r1 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_60_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_59)) begin
                  fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r0 <= in1_din_wire_59;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_60_inst_bnn_fixed_buffer_60_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_59_regbank
         always @(in1_raddr_wire_58 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r0 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r1 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r2 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r3 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r4 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r5 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r6 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r7 or 
fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r8
          or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r9 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r10 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r11 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r12 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r13 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r14 or fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r15)
          begin :fixed_buffer_59_inst
            case (in1_raddr_wire_58) 

               4'd00: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_59_if_1_dout_wire = fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_59_regbank  instance: fixed_buffer_59_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd15) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r15 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd14) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r14 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd13) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r13 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd12) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r12 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd11) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r11 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd10) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r10 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd09) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r9 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd08) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r8 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd07) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r7 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd06) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r6 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd05) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r5 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd04) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r4 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd03) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r3 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd02) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r2 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_58 == 4'd01) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r1 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_59_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_58)) begin
                  fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r0 <= in1_din_wire_58;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_59_inst_bnn_fixed_buffer_59_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_58_regbank
         always @(in1_raddr_wire_57 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r0 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r1 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r2 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r3 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r4 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r5 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r6 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r7 or 
fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r8
          or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r9 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r10 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r11 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r12 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r13 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r14 or fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r15)
          begin :fixed_buffer_58_inst
            case (in1_raddr_wire_57) 

               4'd00: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_58_if_1_dout_wire = fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_58_regbank  instance: fixed_buffer_58_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd15) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r15 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd14) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r14 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd13) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r13 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd12) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r12 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd11) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r11 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd10) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r10 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd09) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r9 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd08) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r8 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd07) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r7 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd06) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r6 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd05) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r5 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd04) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r4 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd03) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r3 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd02) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r2 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_57 == 4'd01) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r1 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_58_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_57)) begin
                  fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r0 <= in1_din_wire_57;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_58_inst_bnn_fixed_buffer_58_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_57_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r0 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r1 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r2 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r3 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r4 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r5 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r6 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r7 or 
fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r8
          or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r9 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r10 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r11 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r12 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r13 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r14 or fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r15)
          begin :fixed_buffer_57_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_57_if_1_dout_wire = fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_57_regbank  instance: fixed_buffer_57_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r15 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r14 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r13 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r12 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r11 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r10 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r9 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r8 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r7 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r6 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r5 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r4 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r3 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r2 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r1 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_57_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r0 <= in1_din_wire_56;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_57_inst_bnn_fixed_buffer_57_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_56_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r0 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r1 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r2 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r3 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r4 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r5 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r6 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r7 or 
fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r8
          or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r9 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r10 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r11 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r12 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r13 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r14 or fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r15)
          begin :fixed_buffer_56_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_56_if_1_dout_wire = fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_56_regbank  instance: fixed_buffer_56_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r15 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r14 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r13 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r12 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r11 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r10 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r9 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r8 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r7 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r6 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r5 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r4 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r3 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r2 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r1 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_56_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r0 <= in1_din_wire_55;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_56_inst_bnn_fixed_buffer_56_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_55_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r0 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r1 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r2 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r3 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r4 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r5 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r6 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r7 or 
fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r8
          or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r9 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r10 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r11 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r12 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r13 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r14 or fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r15)
          begin :fixed_buffer_55_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_55_if_1_dout_wire = fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_55_regbank  instance: fixed_buffer_55_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r15 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r14 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r13 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r12 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r11 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r10 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r9 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r8 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r7 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r6 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r5 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r4 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r3 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r2 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r1 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_55_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r0 <= in1_din_wire_54;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_55_inst_bnn_fixed_buffer_55_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_54_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r0 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r1 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r2 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r3 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r4 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r5 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r6 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r7 or 
fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r8
          or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r9 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r10 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r11 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r12 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r13 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r14 or fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r15)
          begin :fixed_buffer_54_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_54_if_1_dout_wire = fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_54_regbank  instance: fixed_buffer_54_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r15 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r14 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r13 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r12 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r11 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r10 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r9 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r8 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r7 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r6 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r5 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r4 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r3 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r2 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r1 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_54_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r0 <= in1_din_wire_53;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_54_inst_bnn_fixed_buffer_54_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_53_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r0 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r1 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r2 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r3 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r4 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r5 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r6 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r7 or 
fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r8
          or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r9 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r10 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r11 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r12 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r13 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r14 or fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r15)
          begin :fixed_buffer_53_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_53_if_1_dout_wire = fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_53_regbank  instance: fixed_buffer_53_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r15 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r14 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r13 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r12 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r11 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r10 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r9 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r8 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r7 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r6 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r5 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r4 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r3 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r2 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r1 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_53_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r0 <= in1_din_wire_52;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_53_inst_bnn_fixed_buffer_53_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_52_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r0 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r1 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r2 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r3 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r4 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r5 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r6 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r7 or 
fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r8
          or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r9 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r10 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r11 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r12 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r13 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r14 or fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r15)
          begin :fixed_buffer_52_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_52_if_1_dout_wire = fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_52_regbank  instance: fixed_buffer_52_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r15 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r14 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r13 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r12 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r11 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r10 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r9 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r8 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r7 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r6 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r5 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r4 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r3 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r2 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r1 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_52_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r0 <= in1_din_wire_51;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_52_inst_bnn_fixed_buffer_52_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_51_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r0 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r1 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r2 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r3 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r4 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r5 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r6 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r7 or 
fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r8
          or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r9 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r10 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r11 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r12 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r13 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r14 or fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r15)
          begin :fixed_buffer_51_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_51_if_1_dout_wire = fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_51_regbank  instance: fixed_buffer_51_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r15 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r14 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r13 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r12 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r11 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r10 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r9 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r8 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r7 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r6 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r5 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r4 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r3 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r2 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r1 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_51_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r0 <= in1_din_wire_50;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_51_inst_bnn_fixed_buffer_51_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_50_regbank
         always @(in1_raddr_wire_49 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r0 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r1 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r2 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r3 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r4 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r5 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r6 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r7 or 
fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r8
          or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r9 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r10 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r11 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r12 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r13 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r14 or fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r15)
          begin :fixed_buffer_50_inst
            case (in1_raddr_wire_49) 

               4'd00: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_50_if_1_dout_wire = fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_50_regbank  instance: fixed_buffer_50_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd15) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r15 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd14) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r14 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd13) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r13 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd12) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r12 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd11) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r11 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd10) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r10 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd09) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r9 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd08) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r8 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd07) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r7 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd06) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r6 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd05) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r5 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd04) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r4 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd03) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r3 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd02) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r2 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_49 == 4'd01) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r1 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_50_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_49)) begin
                  fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r0 <= in1_din_wire_49;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_50_inst_bnn_fixed_buffer_50_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_49_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r0 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r1 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r2 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r3 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r4 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r5 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r6 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r7 or 
fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r8
          or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r9 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r10 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r11 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r12 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r13 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r14 or fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r15)
          begin :fixed_buffer_49_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_49_if_1_dout_wire = fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_49_regbank  instance: fixed_buffer_49_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r15 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r14 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r13 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r12 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r11 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r10 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r9 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r8 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r7 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r6 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r5 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r4 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r3 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r2 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r1 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_49_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r0 <= in1_din_wire_48;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_49_inst_bnn_fixed_buffer_49_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_48_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r0 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r1 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r2 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r3 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r4 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r5 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r6 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r7 or 
fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r8
          or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r9 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r10 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r11 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r12 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r13 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r14 or fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r15)
          begin :fixed_buffer_48_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_48_if_1_dout_wire = fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_48_regbank  instance: fixed_buffer_48_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r15 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r14 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r13 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r12 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r11 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r10 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r9 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r8 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r7 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r6 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r5 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r4 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r3 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r2 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r1 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_48_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r0 <= in1_din_wire_47;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_48_inst_bnn_fixed_buffer_48_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_47_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r0 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r1 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r2 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r3 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r4 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r5 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r6 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r7 or 
fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r8
          or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r9 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r10 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r11 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r12 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r13 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r14 or fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r15)
          begin :fixed_buffer_47_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_47_if_1_dout_wire = fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_47_regbank  instance: fixed_buffer_47_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r15 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r14 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r13 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r12 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r11 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r10 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r9 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r8 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r7 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r6 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r5 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r4 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r3 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r2 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r1 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_47_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r0 <= in1_din_wire_46;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_47_inst_bnn_fixed_buffer_47_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_46_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r0 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r1 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r2 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r3 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r4 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r5 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r6 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r7 or 
fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r8
          or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r9 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r10 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r11 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r12 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r13 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r14 or fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r15)
          begin :fixed_buffer_46_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_46_if_1_dout_wire = fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_46_regbank  instance: fixed_buffer_46_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r15 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r14 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r13 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r12 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r11 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r10 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r9 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r8 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r7 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r6 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r5 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r4 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r3 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r2 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r1 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_46_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r0 <= in1_din_wire_45;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_46_inst_bnn_fixed_buffer_46_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_45_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r0 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r1 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r2 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r3 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r4 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r5 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r6 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r7 or 
fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r8
          or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r9 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r10 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r11 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r12 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r13 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r14 or fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r15)
          begin :fixed_buffer_45_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_45_if_1_dout_wire = fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_45_regbank  instance: fixed_buffer_45_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r15 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r14 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r13 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r12 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r11 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r10 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r9 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r8 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r7 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r6 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r5 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r4 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r3 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r2 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r1 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_45_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r0 <= in1_din_wire_44;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_45_inst_bnn_fixed_buffer_45_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_44_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r0 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r1 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r2 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r3 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r4 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r5 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r6 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r7 or 
fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r8
          or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r9 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r10 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r11 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r12 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r13 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r14 or fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r15)
          begin :fixed_buffer_44_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_44_if_1_dout_wire = fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_44_regbank  instance: fixed_buffer_44_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r15 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r14 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r13 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r12 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r11 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r10 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r9 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r8 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r7 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r6 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r5 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r4 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r3 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r2 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r1 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_44_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r0 <= in1_din_wire_43;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_44_inst_bnn_fixed_buffer_44_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_43_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r0 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r1 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r2 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r3 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r4 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r5 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r6 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r7 or 
fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r8
          or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r9 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r10 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r11 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r12 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r13 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r14 or fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r15)
          begin :fixed_buffer_43_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_43_if_1_dout_wire = fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_43_regbank  instance: fixed_buffer_43_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r15 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r14 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r13 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r12 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r11 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r10 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r9 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r8 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r7 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r6 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r5 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r4 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r3 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r2 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r1 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_43_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r0 <= in1_din_wire_42;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_43_inst_bnn_fixed_buffer_43_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_42_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r0 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r1 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r2 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r3 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r4 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r5 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r6 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r7 or 
fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r8
          or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r9 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r10 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r11 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r12 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r13 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r14 or fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r15)
          begin :fixed_buffer_42_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_42_if_1_dout_wire = fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_42_regbank  instance: fixed_buffer_42_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r15 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r14 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r13 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r12 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r11 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r10 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r9 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r8 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r7 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r6 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r5 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r4 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r3 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r2 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r1 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_42_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r0 <= in1_din_wire_41;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_42_inst_bnn_fixed_buffer_42_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_41_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r0 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r1 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r2 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r3 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r4 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r5 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r6 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r7 or 
fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r8
          or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r9 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r10 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r11 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r12 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r13 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r14 or fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r15)
          begin :fixed_buffer_41_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_41_if_1_dout_wire = fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_41_regbank  instance: fixed_buffer_41_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r15 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r14 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r13 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r12 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r11 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r10 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r9 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r8 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r7 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r6 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r5 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r4 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r3 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r2 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r1 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_41_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r0 <= in1_din_wire_40;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_41_inst_bnn_fixed_buffer_41_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_40_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r0 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r1 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r2 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r3 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r4 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r5 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r6 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r7 or 
fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r8
          or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r9 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r10 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r11 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r12 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r13 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r14 or fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r15)
          begin :fixed_buffer_40_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_40_if_1_dout_wire = fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_40_regbank  instance: fixed_buffer_40_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r15 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r14 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r13 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r12 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r11 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r10 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r9 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r8 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r7 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r6 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r5 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r4 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r3 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r2 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r1 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_40_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r0 <= in1_din_wire_39;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_40_inst_bnn_fixed_buffer_40_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_39_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r0 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r1 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r2 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r3 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r4 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r5 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r6 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r7 or 
fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r8
          or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r9 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r10 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r11 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r12 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r13 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r14 or fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r15)
          begin :fixed_buffer_39_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_39_if_1_dout_wire = fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_39_regbank  instance: fixed_buffer_39_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r15 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r14 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r13 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r12 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r11 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r10 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r9 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r8 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r7 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r6 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r5 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r4 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r3 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r2 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r1 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_39_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r0 <= in1_din_wire_38;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_39_inst_bnn_fixed_buffer_39_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_38_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r0 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r1 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r2 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r3 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r4 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r5 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r6 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r7 or 
fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r8
          or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r9 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r10 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r11 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r12 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r13 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r14 or fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r15)
          begin :fixed_buffer_38_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_38_if_1_dout_wire = fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_38_regbank  instance: fixed_buffer_38_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r15 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r14 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r13 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r12 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r11 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r10 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r9 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r8 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r7 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r6 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r5 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r4 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r3 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r2 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r1 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_38_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r0 <= in1_din_wire_37;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_38_inst_bnn_fixed_buffer_38_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_37_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r0 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r1 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r2 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r3 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r4 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r5 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r6 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r7 or 
fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r8
          or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r9 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r10 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r11 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r12 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r13 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r14 or fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r15)
          begin :fixed_buffer_37_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_37_if_1_dout_wire = fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_37_regbank  instance: fixed_buffer_37_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r15 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r14 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r13 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r12 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r11 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r10 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r9 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r8 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r7 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r6 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r5 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r4 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r3 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r2 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r1 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_37_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r0 <= in1_din_wire_36;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_37_inst_bnn_fixed_buffer_37_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_36_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r0 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r1 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r2 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r3 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r4 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r5 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r6 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r7 or 
fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r8
          or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r9 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r10 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r11 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r12 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r13 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r14 or fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r15)
          begin :fixed_buffer_36_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_36_if_1_dout_wire = fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_36_regbank  instance: fixed_buffer_36_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r15 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r14 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r13 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r12 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r11 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r10 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r9 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r8 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r7 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r6 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r5 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r4 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r3 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r2 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r1 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_36_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r0 <= in1_din_wire_35;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_36_inst_bnn_fixed_buffer_36_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_35_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r0 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r1 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r2 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r3 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r4 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r5 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r6 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r7 or 
fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r8
          or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r9 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r10 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r11 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r12 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r13 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r14 or fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r15)
          begin :fixed_buffer_35_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_35_if_1_dout_wire = fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_35_regbank  instance: fixed_buffer_35_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r15 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r14 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r13 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r12 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r11 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r10 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r9 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r8 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r7 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r6 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r5 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r4 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r3 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r2 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r1 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_35_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r0 <= in1_din_wire_34;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_35_inst_bnn_fixed_buffer_35_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_34_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r0 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r1 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r2 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r3 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r4 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r5 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r6 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r7 or 
fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r8
          or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r9 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r10 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r11 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r12 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r13 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r14 or fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r15)
          begin :fixed_buffer_34_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_34_if_1_dout_wire = fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_34_regbank  instance: fixed_buffer_34_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r15 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r14 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r13 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r12 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r11 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r10 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r9 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r8 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r7 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r6 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r5 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r4 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r3 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r2 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r1 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_34_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r0 <= in1_din_wire_33;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_34_inst_bnn_fixed_buffer_34_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_33_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r0 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r1 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r2 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r3 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r4 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r5 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r6 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r7 or 
fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r8
          or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r9 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r10 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r11 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r12 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r13 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r14 or fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r15)
          begin :fixed_buffer_33_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_33_if_1_dout_wire = fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_33_regbank  instance: fixed_buffer_33_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r15 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r14 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r13 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r12 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r11 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r10 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r9 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r8 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r7 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r6 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r5 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r4 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r3 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r2 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r1 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_33_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r0 <= in1_din_wire_32;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_33_inst_bnn_fixed_buffer_33_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_32_regbank
         always @(in1_raddr_wire_31 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r0 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r1 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r2 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r3 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r4 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r5 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r6 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r7 or 
fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r8
          or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r9 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r10 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r11 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r12 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r13 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r14 or fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r15)
          begin :fixed_buffer_32_inst
            case (in1_raddr_wire_31) 

               4'd00: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_32_if_1_dout_wire = fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_32_regbank  instance: fixed_buffer_32_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd15) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r15 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd14) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r14 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd13) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r13 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd12) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r12 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd11) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r11 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd10) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r10 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd09) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r9 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd08) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r8 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd07) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r7 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd06) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r6 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd05) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r5 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd04) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r4 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd03) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r3 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd02) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r2 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && in2_waddr_wire_31 == 4'd01) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r1 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_32_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_32_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire_31)) begin
                  fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r0 <= in1_din_wire_31;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_32_inst_bnn_fixed_buffer_32_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_31_regbank
         always @(in1_raddr_wire or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r0 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r1 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r2 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r3 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r4 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r5 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r6 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r7 or 
fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r8
          or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r9 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r10 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r11 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r12 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r13 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r14 or fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r15)
          begin :fixed_buffer_31_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_31_if_1_dout_wire = fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_31_regbank  instance: fixed_buffer_31_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r15 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r14 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r13 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r12 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r11 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r10 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r9 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r8 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r7 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r6 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r5 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r4 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r3 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r2 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r1 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_31_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r0 <= in1_din_wire_30;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_31_inst_bnn_fixed_buffer_31_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_30_regbank
         always @(in1_raddr_wire or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r0 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r1 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r2 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r3 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r4 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r5 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r6 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r7 or 
fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r8
          or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r9 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r10 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r11 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r12 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r13 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r14 or fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r15)
          begin :fixed_buffer_30_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_30_if_1_dout_wire = fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_30_regbank  instance: fixed_buffer_30_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r15 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r14 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r13 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r12 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r11 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r10 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r9 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r8 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r7 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r6 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r5 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r4 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r3 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r2 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r1 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_30_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r0 <= in1_din_wire_29;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_30_inst_bnn_fixed_buffer_30_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_29_regbank
         always @(in1_raddr_wire or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r0 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r1 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r2 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r3 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r4 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r5 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r6 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r7 or 
fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r8
          or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r9 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r10 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r11 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r12 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r13 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r14 or fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r15)
          begin :fixed_buffer_29_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_29_if_1_dout_wire = fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_29_regbank  instance: fixed_buffer_29_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r15 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r14 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r13 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r12 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r11 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r10 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r9 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r8 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r7 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r6 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r5 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r4 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r3 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r2 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r1 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_29_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r0 <= in1_din_wire_28;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_29_inst_bnn_fixed_buffer_29_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_28_regbank
         always @(in1_raddr_wire or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r0 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r1 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r2 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r3 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r4 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r5 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r6 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r7 or 
fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r8
          or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r9 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r10 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r11 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r12 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r13 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r14 or fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r15)
          begin :fixed_buffer_28_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_28_if_1_dout_wire = fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_28_regbank  instance: fixed_buffer_28_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r15 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r14 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r13 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r12 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r11 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r10 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r9 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r8 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r7 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r6 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r5 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r4 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r3 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r2 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r1 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_28_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r0 <= in1_din_wire_27;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_28_inst_bnn_fixed_buffer_28_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_27_regbank
         always @(in1_raddr_wire or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r0 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r1 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r2 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r3 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r4 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r5 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r6 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r7 or 
fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r8
          or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r9 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r10 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r11 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r12 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r13 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r14 or fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r15)
          begin :fixed_buffer_27_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_27_if_1_dout_wire = fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_27_regbank  instance: fixed_buffer_27_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r15 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r14 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r13 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r12 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r11 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r10 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r9 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r8 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r7 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r6 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r5 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r4 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r3 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r2 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r1 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_27_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r0 <= in1_din_wire_26;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_27_inst_bnn_fixed_buffer_27_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_26_regbank
         always @(in1_raddr_wire or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r0 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r1 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r2 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r3 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r4 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r5 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r6 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r7 or 
fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r8
          or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r9 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r10 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r11 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r12 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r13 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r14 or fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r15)
          begin :fixed_buffer_26_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_26_if_1_dout_wire = fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_26_regbank  instance: fixed_buffer_26_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r15 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r14 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r13 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r12 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r11 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r10 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r9 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r8 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r7 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r6 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r5 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r4 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r3 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r2 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r1 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_26_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r0 <= in1_din_wire_25;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_26_inst_bnn_fixed_buffer_26_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_25_regbank
         always @(in1_raddr_wire or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r0 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r1 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r2 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r3 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r4 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r5 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r6 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r7 or 
fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r8
          or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r9 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r10 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r11 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r12 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r13 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r14 or fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r15)
          begin :fixed_buffer_25_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_25_if_1_dout_wire = fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_25_regbank  instance: fixed_buffer_25_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r15 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r14 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r13 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r12 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r11 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r10 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r9 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r8 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r7 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r6 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r5 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r4 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r3 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r2 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r1 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_25_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r0 <= in1_din_wire_24;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_25_inst_bnn_fixed_buffer_25_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_24_regbank
         always @(in1_raddr_wire or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r0 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r1 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r2 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r3 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r4 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r5 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r6 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r7 or 
fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r8
          or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r9 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r10 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r11 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r12 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r13 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r14 or fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r15)
          begin :fixed_buffer_24_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_24_if_1_dout_wire = fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_24_regbank  instance: fixed_buffer_24_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r15 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r14 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r13 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r12 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r11 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r10 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r9 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r8 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r7 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r6 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r5 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r4 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r3 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r2 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r1 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_24_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r0 <= in1_din_wire_23;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_24_inst_bnn_fixed_buffer_24_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_23_regbank
         always @(in1_raddr_wire or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r0 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r1 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r2 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r3 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r4 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r5 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r6 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r7 or 
fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r8
          or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r9 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r10 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r11 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r12 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r13 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r14 or fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r15)
          begin :fixed_buffer_23_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_23_if_1_dout_wire = fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_23_regbank  instance: fixed_buffer_23_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r15 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r14 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r13 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r12 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r11 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r10 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r9 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r8 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r7 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r6 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r5 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r4 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r3 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r2 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r1 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_23_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r0 <= in1_din_wire_22;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_23_inst_bnn_fixed_buffer_23_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_22_regbank
         always @(in1_raddr_wire or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r0 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r1 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r2 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r3 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r4 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r5 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r6 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r7 or 
fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r8
          or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r9 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r10 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r11 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r12 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r13 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r14 or fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r15)
          begin :fixed_buffer_22_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_22_if_1_dout_wire = fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_22_regbank  instance: fixed_buffer_22_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r15 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r14 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r13 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r12 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r11 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r10 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r9 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r8 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r7 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r6 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r5 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r4 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r3 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r2 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r1 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_22_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r0 <= in1_din_wire_21;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_22_inst_bnn_fixed_buffer_22_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_21_regbank
         always @(in1_raddr_wire or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r0 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r1 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r2 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r3 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r4 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r5 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r6 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r7 or 
fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r8
          or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r9 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r10 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r11 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r12 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r13 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r14 or fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r15)
          begin :fixed_buffer_21_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_21_if_1_dout_wire = fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_21_regbank  instance: fixed_buffer_21_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r15 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r14 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r13 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r12 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r11 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r10 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r9 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r8 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r7 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r6 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r5 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r4 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r3 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r2 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r1 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_21_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r0 <= in1_din_wire_20;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_21_inst_bnn_fixed_buffer_21_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_20_regbank
         always @(in1_raddr_wire or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r0 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r1 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r2 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r3 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r4 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r5 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r6 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r7 or 
fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r8
          or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r9 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r10 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r11 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r12 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r13 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r14 or fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r15)
          begin :fixed_buffer_20_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_20_if_1_dout_wire = fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_20_regbank  instance: fixed_buffer_20_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r15 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r14 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r13 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r12 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r11 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r10 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r9 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r8 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r7 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r6 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r5 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r4 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r3 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r2 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r1 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_20_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r0 <= in1_din_wire_19;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_20_inst_bnn_fixed_buffer_20_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_19_regbank
         always @(in1_raddr_wire or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r0 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r1 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r2 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r3 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r4 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r5 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r6 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r7 or 
fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r8
          or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r9 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r10 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r11 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r12 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r13 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r14 or fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r15)
          begin :fixed_buffer_19_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_19_if_1_dout_wire = fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_19_regbank  instance: fixed_buffer_19_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r15 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r14 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r13 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r12 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r11 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r10 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r9 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r8 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r7 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r6 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r5 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r4 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r3 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r2 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r1 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_19_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r0 <= in1_din_wire_18;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_19_inst_bnn_fixed_buffer_19_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_18_regbank
         always @(in1_raddr_wire or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r0 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r1 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r2 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r3 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r4 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r5 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r6 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r7 or 
fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r8
          or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r9 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r10 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r11 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r12 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r13 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r14 or fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r15)
          begin :fixed_buffer_18_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_18_if_1_dout_wire = fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_18_regbank  instance: fixed_buffer_18_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r15 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r14 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r13 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r12 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r11 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r10 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r9 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r8 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r7 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r6 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r5 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r4 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r3 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r2 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r1 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_18_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r0 <= in1_din_wire_17;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_18_inst_bnn_fixed_buffer_18_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_17_regbank
         always @(in1_raddr_wire or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r0 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r1 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r2 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r3 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r4 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r5 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r6 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r7 or 
fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r8
          or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r9 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r10 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r11 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r12 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r13 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r14 or fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r15)
          begin :fixed_buffer_17_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_17_if_1_dout_wire = fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_17_regbank  instance: fixed_buffer_17_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r15 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r14 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r13 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r12 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r11 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r10 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r9 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r8 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r7 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r6 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r5 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r4 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r3 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r2 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r1 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_17_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r0 <= in1_din_wire_16;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_17_inst_bnn_fixed_buffer_17_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_16_regbank
         always @(in1_raddr_wire or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r0 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r1 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r2 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r3 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r4 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r5 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r6 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r7 or 
fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r8
          or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r9 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r10 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r11 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r12 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r13 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r14 or fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r15)
          begin :fixed_buffer_16_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_16_if_1_dout_wire = fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_16_regbank  instance: fixed_buffer_16_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r15 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r14 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r13 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r12 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r11 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r10 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r9 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r8 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r7 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r6 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r5 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r4 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r3 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r2 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r1 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_16_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r0 <= in1_din_wire_15;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_16_inst_bnn_fixed_buffer_16_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_15_regbank
         always @(in1_raddr_wire or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r0 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r1 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r2 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r3 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r4 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r5 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r6 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r7 or 
fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r8
          or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r9 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r10 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r11 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r12 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r13 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r14 or fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r15)
          begin :fixed_buffer_15_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_15_if_1_dout_wire = fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_15_regbank  instance: fixed_buffer_15_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r15 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r14 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r13 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r12 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r11 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r10 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r9 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r8 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r7 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r6 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r5 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r4 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r3 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r2 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r1 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_15_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r0 <= in1_din_wire_14;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_15_inst_bnn_fixed_buffer_15_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_14_regbank
         always @(in1_raddr_wire or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r0 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r1 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r2 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r3 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r4 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r5 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r6 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r7 or 
fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r8
          or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r9 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r10 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r11 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r12 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r13 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r14 or fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r15)
          begin :fixed_buffer_14_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_14_if_1_dout_wire = fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_14_regbank  instance: fixed_buffer_14_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r15 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r14 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r13 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r12 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r11 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r10 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r9 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r8 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r7 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r6 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r5 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r4 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r3 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r2 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r1 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_14_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r0 <= in1_din_wire_13;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_14_inst_bnn_fixed_buffer_14_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_13_regbank
         always @(in1_raddr_wire or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r0 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r1 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r2 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r3 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r4 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r5 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r6 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r7 or 
fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r8
          or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r9 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r10 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r11 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r12 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r13 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r14 or fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r15)
          begin :fixed_buffer_13_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_13_if_1_dout_wire = fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_13_regbank  instance: fixed_buffer_13_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r15 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r14 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r13 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r12 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r11 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r10 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r9 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r8 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r7 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r6 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r5 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r4 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r3 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r2 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r1 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_13_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r0 <= in1_din_wire_12;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_13_inst_bnn_fixed_buffer_13_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_12_regbank
         always @(in1_raddr_wire or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r0 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r1 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r2 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r3 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r4 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r5 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r6 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r7 or 
fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r8
          or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r9 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r10 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r11 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r12 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r13 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r14 or fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r15)
          begin :fixed_buffer_12_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_12_if_1_dout_wire = fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_12_regbank  instance: fixed_buffer_12_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r15 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r14 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r13 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r12 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r11 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r10 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r9 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r8 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r7 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r6 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r5 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r4 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r3 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r2 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r1 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_12_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r0 <= in1_din_wire_11;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_12_inst_bnn_fixed_buffer_12_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_11_regbank
         always @(in1_raddr_wire or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r0 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r1 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r2 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r3 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r4 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r5 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r6 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r7 or 
fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r8
          or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r9 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r10 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r11 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r12 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r13 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r14 or fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r15)
          begin :fixed_buffer_11_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_11_if_1_dout_wire = fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_11_regbank  instance: fixed_buffer_11_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r15 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r14 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r13 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r12 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r11 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r10 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r9 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r8 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r7 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r6 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r5 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r4 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r3 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r2 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r1 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_11_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r0 <= in1_din_wire_10;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_11_inst_bnn_fixed_buffer_11_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_10_regbank
         always @(in1_raddr_wire or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r0 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r1 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r2 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r3 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r4 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r5 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r6 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r7 or 
fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r8
          or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r9 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r10 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r11 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r12 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r13 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r14 or fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r15)
          begin :fixed_buffer_10_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_10_if_1_dout_wire = fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_10_regbank  instance: fixed_buffer_10_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r15 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r14 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r13 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r12 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r11 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r10 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r9 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r8 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r7 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r6 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r5 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r4 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r3 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r2 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r1 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_10_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r0 <= in1_din_wire_9;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_10_inst_bnn_fixed_buffer_10_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_9_regbank
         always @(in1_raddr_wire or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r0 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r1 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r2 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r3 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r4 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r5 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r6 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r7 or 
fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r8
          or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r9 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r10 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r11 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r12 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r13 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r14 or fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r15)
          begin :fixed_buffer_9_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_9_if_1_dout_wire = fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_9_regbank  instance: fixed_buffer_9_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r15 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r14 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r13 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r12 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r11 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r10 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r9 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r8 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r7 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r6 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r5 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r4 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r3 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r2 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r1 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_9_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r0 <= in1_din_wire_8;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_9_inst_bnn_fixed_buffer_9_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_8_regbank
         always @(in1_raddr_wire or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r0 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r1 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r2 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r3 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r4 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r5 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r6 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r7 or 
fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r8
          or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r9 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r10 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r11 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r12 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r13 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r14 or fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r15)
          begin :fixed_buffer_8_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_8_if_1_dout_wire = fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_8_regbank  instance: fixed_buffer_8_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r15 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r14 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r13 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r12 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r11 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r10 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r9 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r8 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r7 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r6 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r5 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r4 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r3 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r2 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r1 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_8_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r0 <= in1_din_wire_7;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_8_inst_bnn_fixed_buffer_8_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_7_regbank
         always @(in1_raddr_wire or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r0 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r1 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r2 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r3 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r4 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r5 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r6 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r7 or 
fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r8
          or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r9 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r10 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r11 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r12 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r13 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r14 or fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r15)
          begin :fixed_buffer_7_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_7_if_1_dout_wire = fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_7_regbank  instance: fixed_buffer_7_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r15 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r14 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r13 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r12 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r11 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r10 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r9 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r8 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r7 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r6 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r5 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r4 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r3 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r2 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r1 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_7_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r0 <= in1_din_wire_6;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_7_inst_bnn_fixed_buffer_7_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_6_regbank
         always @(in1_raddr_wire or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r0 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r1 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r2 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r3 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r4 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r5 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r6 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r7 or 
fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r8
          or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r9 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r10 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r11 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r12 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r13 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r14 or fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r15)
          begin :fixed_buffer_6_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_6_if_1_dout_wire = fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_6_regbank  instance: fixed_buffer_6_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r15 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r14 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r13 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r12 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r11 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r10 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r9 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r8 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r7 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r6 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r5 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r4 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r3 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r2 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r1 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_6_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r0 <= in1_din_wire_5;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_6_inst_bnn_fixed_buffer_6_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_5_regbank
         always @(in1_raddr_wire or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r0 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r1 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r2 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r3 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r4 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r5 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r6 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r7 or 
fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r8
          or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r9 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r10 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r11 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r12 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r13 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r14 or fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r15)
          begin :fixed_buffer_5_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_5_if_1_dout_wire = fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_5_regbank  instance: fixed_buffer_5_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r15 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r14 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r13 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r12 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r11 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r10 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r9 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r8 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r7 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r6 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r5 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r4 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r3 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r2 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r1 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_5_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r0 <= in1_din_wire_4;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_5_inst_bnn_fixed_buffer_5_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_4_regbank
         always @(in1_raddr_wire or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r0 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r1 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r2 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r3 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r4 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r5 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r6 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r7 or 
fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r8
          or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r9 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r10 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r11 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r12 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r13 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r14 or fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r15)
          begin :fixed_buffer_4_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_4_if_1_dout_wire = fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_4_regbank  instance: fixed_buffer_4_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r15 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r14 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r13 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r12 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r11 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r10 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r9 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r8 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r7 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r6 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r5 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r4 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r3 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r2 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r1 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_4_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r0 <= in1_din_wire_3;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_4_inst_bnn_fixed_buffer_4_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_3_regbank
         always @(in1_raddr_wire or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r0 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r1 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r2 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r3 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r4 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r5 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r6 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r7 or 
fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r8
          or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r9 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r10 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r11 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r12 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r13 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r14 or fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r15)
          begin :fixed_buffer_3_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_3_if_1_dout_wire = fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_3_regbank  instance: fixed_buffer_3_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r15 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r14 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r13 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r12 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r11 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r10 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r9 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r8 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r7 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r6 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r5 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r4 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r3 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r2 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r1 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_3_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r0 <= in1_din_wire_2;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_3_inst_bnn_fixed_buffer_3_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_2_regbank
         always @(in1_raddr_wire or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r0 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r1 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r2 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r3 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r4 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r5 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r6 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r7 or 
fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r8
          or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r9 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r10 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r11 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r12 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r13 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r14 or fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r15)
          begin :fixed_buffer_2_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_2_if_1_dout_wire = fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_2_regbank  instance: fixed_buffer_2_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r15 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r14 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r13 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r12 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r11 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r10 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r9 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r8 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r7 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r6 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r5 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r4 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r3 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r2 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r1 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_2_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r0 <= in1_din_wire_1;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_2_inst_bnn_fixed_buffer_2_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_1_regbank
         always @(in1_raddr_wire or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r0 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r1 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r2 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r3 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r4 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r5 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r6 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r7 or 
fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r8
          or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r9 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r10 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r11 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r12 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r13 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r14 or fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r15)
          begin :fixed_buffer_1_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_1_if_1_dout_wire = fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_1_regbank  instance: fixed_buffer_1_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r15 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r14 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r13 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r12 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r11 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r10 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r9 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r8 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r7 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r6 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r5 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r4 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r3 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r2 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r1 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_1_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r0 <= in1_din_wire_0;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_1_inst_bnn_fixed_buffer_1_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         // resource: bnn_fixed_buffer_0_regbank
         always @(in1_raddr_wire or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r0 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r1 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r2 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r3 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r4 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r5 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r6 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r7 or 
fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r8
          or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r9 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r10 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r11 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r12 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r13 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r14 or fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r15)
          begin :fixed_buffer_0_inst
            case (in1_raddr_wire) 

               4'd00: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r0;
               end
               
               4'd01: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r1;
               end
               
               4'd02: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r2;
               end
               
               4'd03: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r3;
               end
               
               4'd04: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r4;
               end
               
               4'd05: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r5;
               end
               
               4'd06: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r6;
               end
               
               4'd07: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r7;
               end
               
               4'd08: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r8;
               end
               
               4'd09: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r9;
               end
               
               4'd10: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r10;
               end
               
               4'd11: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r11;
               end
               
               4'd12: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r12;
               end
               
               4'd13: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r13;
               end
               
               4'd14: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r14;
               end
               
               4'd15: begin
                  fixed_buffer_0_if_1_dout_wire = fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r15;
               end
               
            endcase

         end

         // resource: bnn_fixed_buffer_0_regbank  instance: fixed_buffer_0_inst
         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r15
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd15) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r15 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd15) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r15 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r14
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd14) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r14 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd14) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r14 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r13
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd13) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r13 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd13) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r13 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r12
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd12) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r12 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd12) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r12 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r11
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd11) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r11 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd11) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r11 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r10
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd10) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r10 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd10) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r10 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r9
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd09) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r9 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd09) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r9 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r8
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd08) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r8 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd08) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r8 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r7
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd07) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r7 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd07) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r7 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r6
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd06) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r6 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd06) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r6 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r5
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd05) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r5 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd05) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r5 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r4
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd04) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r4 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd04) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r4 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r3
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd03) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r3 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd03) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r3 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r2
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd02) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r2 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd02) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r2 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r1
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && in2_waddr_wire == 4'd01) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r1 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && in1_waddr_wire == 4'd01) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r1 <= 12'd0000;
                  end
               end
            end
         end

         always @(posedge clk)
          begin :write_bnn_fixed_buffer_0_regbank_r0
            if (stall0) begin
            end
            else begin
               if (fixed_buffer_0_if_2_wen0_wire == 1'b1 && !(|in2_waddr_wire)) begin
                  fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r0 <= in1_din_wire;
               end
               else begin
                  if (fixed_buffer_0_if_0_wen0_wire == 1'b1 && !(|in1_waddr_wire)) begin
                     fixed_buffer_0_inst_bnn_fixed_buffer_0_regbank_r0 <= 12'd0000;
                  end
               end
            end
         end

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5019(
                               .in2( bnn_Mod_6Ux32U_7U_4_5019_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5019_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5018(
                               .in2( bnn_Mod_6Ux32U_7U_4_5018_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5018_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5017(
                               .in2( bnn_Mod_6Ux32U_7U_4_5017_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5017_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5016(
                               .in2( bnn_Mod_6Ux32U_7U_4_5016_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5016_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5015(
                               .in2( bnn_Mod_6Ux32U_7U_4_5015_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5015_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5014(
                               .in2( bnn_Mod_6Ux32U_7U_4_5014_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5014_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5013(
                               .in2( bnn_Mod_6Ux32U_7U_4_5013_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5013_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5012(
                               .in2( bnn_Mod_6Ux32U_7U_4_5012_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5012_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5011(
                               .in2( bnn_Mod_6Ux32U_7U_4_5011_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5011_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5010(
                               .in2( bnn_Mod_6Ux32U_7U_4_5010_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5010_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5009(
                               .in2( bnn_Mod_6Ux32U_7U_4_5009_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5009_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5008(
                               .in2( bnn_Mod_6Ux32U_7U_4_5008_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5008_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5007(
                               .in2( bnn_Mod_6Ux32U_7U_4_5007_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5007_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5006(
                               .in2( bnn_Mod_6Ux32U_7U_4_5006_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5006_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5005(
                               .in2( bnn_Mod_6Ux32U_7U_4_5005_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5005_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5004(
                               .in2( bnn_Mod_6Ux32U_7U_4_5004_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5004_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5003(
                               .in2( bnn_Mod_6Ux32U_7U_4_5003_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5003_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5002(
                               .in2( bnn_Mod_6Ux32U_7U_4_5002_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5002_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5001(
                               .in2( bnn_Mod_6Ux32U_7U_4_5001_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5001_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_5000(
                               .in2( bnn_Mod_6Ux32U_7U_4_5000_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_5000_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4999(
                               .in2( bnn_Mod_6Ux32U_7U_4_4999_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4999_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4998(
                               .in2( bnn_Mod_6Ux32U_7U_4_4998_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4998_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4997(
                               .in2( bnn_Mod_6Ux32U_7U_4_4997_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4997_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4996(
                               .in2( bnn_Mod_6Ux32U_7U_4_4996_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4996_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4995(
                               .in2( bnn_Mod_6Ux32U_7U_4_4995_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4995_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4994(
                               .in2( bnn_Mod_6Ux32U_7U_4_4994_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4994_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4993(
                               .in2( bnn_Mod_6Ux32U_7U_4_4993_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4993_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4992(
                               .in2( bnn_Mod_6Ux32U_7U_4_4992_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4992_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4991(
                               .in2( bnn_Mod_6Ux32U_7U_4_4991_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4991_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4990(
                               .in2( bnn_Mod_6Ux32U_7U_4_4990_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4990_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4989(
                               .in2( bnn_Mod_6Ux32U_7U_4_4989_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4989_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         bnn_Mod_6Ux32U_7U_4 bnn_Mod_6Ux32U_7U_4_4988(
                               .in2( bnn_Mod_6Ux32U_7U_4_4988_in2 ),
                               .in1( s_reg_1002 ),
                               .out1( bnn_Mod_6Ux32U_7U_4_4988_out1 ),
                               .clk( clk ),
                               .stall( stall0 )
                             );

         
// pragma translate_off
         always @(posedge clk)
          begin :drive_printf
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_GreaterThan_32Ux6U_1U_4_179_out1) begin
                        $write("%s:%d: assertion failure\n", "bnn.cc", 9'd164);
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        $write("==== Finished Accel ====\n");
                     end
                  end
                  
                  5'd19: begin
                     if (en_2) begin
                        case (cycle2_state2) 

                           2'd0, 2'd1: begin
                              if (s_reg_870_stage10) begin
                              end
                              else begin
                                 $write("===== Entering Accel =====\n");
                                 if (bnn_GreaterThan_64Ux10U_1U_4_149_out1) begin
                                    $write("%s:%d: assertion failure\n", "bnn.cc", 9'd162);
                                 end
                              end
                           end
                           
                        endcase

                     end
                  end
                  
               endcase

            end
         end
// pragma translate_on

         // resource: mux_97bx8i
         // resource: regr_97b
         always @(posedge clk)
          begin :drive_memreq_data
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     memreq_data_slice <= {{1'b0, s_reg_1007}, 64'd00000000000000000000};
                  end
                  
                  5'd02: begin
                     memreq_data_slice <= {{1'b0, s_reg_1017}, 64'd00000000000000000000};
                  end
                  
                  5'd04: begin
                     memreq_data_slice <= {{1'b0, s_reg_1008}, 64'd00000000000000000000};
                  end
                  
                  5'd11: begin
                     memreq_data_slice <= {{1'b0, bnn_Add_32Ux32U_32U_1_955_out1}, 64'd00000000000000000000};
                  end
                  
                  5'd12: begin
                     if (bnn_LessThan_10Ux32U_1U_4_4104_out1) begin
                        memreq_data_slice <= {{1'b0, bnn_Add_32Ux10U_32U_1_954_out1}, 64'd00000000000000000000};
                     end
                     else begin
                        memreq_data_slice <= {{1'b0, s_reg_1008}, 64'd00000000000000000000};
                     end
                  end
                  
                  5'd14, 5'd18: begin
                     memreq_data_slice <= {1'b1, {bnn_Add_32Ux32U_32U_1_955_out1, {{ 52 {bnn_N_Mux_12_64_13_4_5206_out1[11]}}, bnn_N_Mux_12_64_13_4_5206_out1}}};
                  end
                  
                  5'd15: begin
                     if (!cycle3_state && !s_reg_1044_stage2) begin
                        memreq_data_slice <= {1'b1, {bnn_Add_32Ux32U_32U_1_955_out1, {{ 52 {bnn_N_Mux_12_64_13_4_5206_out1[11]}}, bnn_N_Mux_12_64_13_4_5206_out1}}};
                     end
                     else begin
                        memreq_data_slice <= {1'b1, {s_reg_1001, bnn_And_64Sx64S_64S_1_5201_out1}};
                     end
                  end
                  
                  5'd16: begin
                     if (!cycle2_state1 && !s_reg_907) begin
                        if (drain) begin
                           memreq_data_slice <= {1'b1, {bnn_Add_32Ux32U_32U_1_955_out1, {{ 52 {bnn_N_Mux_12_64_13_4_5206_out1[11]}}, bnn_N_Mux_12_64_13_4_5206_out1}}};
                        end
                        else begin
                           memreq_data_slice <= {1'b1, {bnn_Add_32Ux10U_32U_1_954_out1, {bnn_Add_17Sx16S_17S_1_3146_out1[16], {bnn_Add_17Sx16S_17S_1_3128_out1[16], {bnn_Add_17Sx16S_17S_1_3107_out1[16], {bnn_Add_17Sx16S_17S_1_3083_out1[16], {bnn_Add_17Sx16S_17S_1_3057_out1[16], {bnn_Add_17Sx16S_17S_1_3030_out1[16], {bnn_Add_17Sx16S_17S_1_3005_out1[16], {bnn_Add_17Sx16S_17S_1_2981_out1[16], {bnn_Add_17Sx16S_17S_1_2957_out1[16], {bnn_Add_17Sx16S_17S_1_2932_out1[16], {bnn_Add_17Sx16S_17S_1_2905_out1
[
                           16], {bnn_Add_17Sx16S_17S_1_2878_out1[16], {bnn_Add_17Sx16S_17S_1_2851_out1[16], {bnn_Add_17Sx16S_17S_1_2824_out1[16], {bnn_Add_17Sx16S_17S_1_2797_out1[16], {bnn_Add_17Sx16S_17S_1_2769_out1[16], {bnn_Add_17Sx16S_17S_1_2741_out1[16], {bnn_Add_17Sx16S_17S_1_2714_out1[16], {bnn_Add_17Sx16S_17S_1_2687_out1[16], {bnn_Add_17Sx16S_17S_1_2660_out1[16], {bnn_Add_17Sx16S_17S_1_2633_out1[16], {bnn_Add_17Sx16S_17S_1_2606_out1[16], {bnn_Add_17Sx16S_17S_1_2579_out1[16]
                               , {bnn_Add_17Sx16S_17S_1_2552_out1[16], {bnn_Add_17Sx16S_17S_1_2525_out1[16], {bnn_Add_17Sx16S_17S_1_2498_out1[16], {bnn_Add_17Sx16S_17S_1_2471_out1[16], {bnn_Add_17Sx16S_17S_1_2444_out1[16], {bnn_Add_17Sx16S_17S_1_2417_out1[16], {bnn_Add_17Sx16S_17S_1_2390_out1[16], {bnn_Add_17Sx16S_17S_1_3547_out1[16], {bnn_Add_17Sx16S_17S_1_3546_out1[16], {bnn_Add_17Sx16S_17S_1_3542_out1[16], {bnn_Add_17Sx16S_17S_1_3534_out1[16], {bnn_Add_17Sx16S_17S_1_3521_out1[16]
                               , {bnn_Add_17Sx16S_17S_1_3506_out1[16], {bnn_Add_17Sx16S_17S_1_3491_out1[16], {bnn_Add_17Sx16S_17S_1_3477_out1[16], {bnn_Add_17Sx16S_17S_1_3464_out1[16], {bnn_Add_17Sx16S_17S_1_3451_out1[16], {bnn_Add_17Sx16S_17S_1_3436_out1[16], {bnn_Add_17Sx16S_17S_1_3418_out1[16], {bnn_Add_17Sx16S_17S_1_3400_out1[16], {bnn_Add_17Sx16S_17S_1_3384_out1[16], {bnn_Add_17Sx16S_17S_1_3369_out1[16], {bnn_Add_17Sx16S_17S_1_3355_out1[16], {bnn_Add_17Sx16S_17S_1_3342_out1[16]
                               , {bnn_Add_17Sx16S_17S_1_3329_out1[16], {bnn_Add_17Sx16S_17S_1_3233_out1[16], {bnn_Add_17Sx16S_17S_1_3220_out1[16], {bnn_Add_17Sx16S_17S_1_3207_out1[16], {bnn_Add_17Sx16S_17S_1_3192_out1[16], {bnn_Add_17Sx16S_17S_1_3174_out1[16], {bnn_Add_17Sx16S_17S_1_3155_out1[16], {bnn_Add_17Sx16S_17S_1_3137_out1[16], {bnn_Add_17Sx16S_17S_1_3097_out1[16], {bnn_Add_17Sx16S_17S_1_3296_out1[16], {bnn_Add_17Sx16S_17S_1_3262_out1[16], {bnn_Add_17Sx16S_17S_1_3247_out1[16]
                               , {bnn_Add_17Sx16S_17S_1_3278_out1[16], {bnn_Add_17Sx16S_17S_1_3314_out1[16], {bnn_Add_17Sx16S_17S_1_3118_out1[16], {bnn_Add_17Sx16S_17S_1_3162_out1[16], bnn_Add_17Sx16S_17S_1_2389_out1[16]}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}};
                        end
                     end
                     else begin
                        memreq_data_slice <= {1'b1, {bnn_Add_32Ux10U_32U_1_954_out1, {bnn_Add_17Sx16S_17S_1_3146_out1[16], {bnn_Add_17Sx16S_17S_1_3128_out1[16], {bnn_Add_17Sx16S_17S_1_3107_out1[16], {bnn_Add_17Sx16S_17S_1_3083_out1[16], {bnn_Add_17Sx16S_17S_1_3057_out1[16], {bnn_Add_17Sx16S_17S_1_3030_out1[16], {bnn_Add_17Sx16S_17S_1_3005_out1[16], {bnn_Add_17Sx16S_17S_1_2981_out1[16], {bnn_Add_17Sx16S_17S_1_2957_out1[16], {bnn_Add_17Sx16S_17S_1_2932_out1[16], {bnn_Add_17Sx16S_17S_1_2905_out1
                            [16], {bnn_Add_17Sx16S_17S_1_2878_out1[16], {bnn_Add_17Sx16S_17S_1_2851_out1[16], {bnn_Add_17Sx16S_17S_1_2824_out1[16], {bnn_Add_17Sx16S_17S_1_2797_out1[16], {bnn_Add_17Sx16S_17S_1_2769_out1[16], {bnn_Add_17Sx16S_17S_1_2741_out1[16], {bnn_Add_17Sx16S_17S_1_2714_out1[16], {bnn_Add_17Sx16S_17S_1_2687_out1[16], {bnn_Add_17Sx16S_17S_1_2660_out1[16], {bnn_Add_17Sx16S_17S_1_2633_out1[16], {bnn_Add_17Sx16S_17S_1_2606_out1[16], {bnn_Add_17Sx16S_17S_1_2579_out1[16]
                            , {bnn_Add_17Sx16S_17S_1_2552_out1[16], {bnn_Add_17Sx16S_17S_1_2525_out1[16], {bnn_Add_17Sx16S_17S_1_2498_out1[16], {bnn_Add_17Sx16S_17S_1_2471_out1[16], {bnn_Add_17Sx16S_17S_1_2444_out1[16], {bnn_Add_17Sx16S_17S_1_2417_out1[16], {bnn_Add_17Sx16S_17S_1_2390_out1[16], {bnn_Add_17Sx16S_17S_1_3547_out1[16], {bnn_Add_17Sx16S_17S_1_3546_out1[16], {bnn_Add_17Sx16S_17S_1_3542_out1[16], {bnn_Add_17Sx16S_17S_1_3534_out1[16], {bnn_Add_17Sx16S_17S_1_3521_out1[16]
                            , {bnn_Add_17Sx16S_17S_1_3506_out1[16], {bnn_Add_17Sx16S_17S_1_3491_out1[16], {bnn_Add_17Sx16S_17S_1_3477_out1[16], {bnn_Add_17Sx16S_17S_1_3464_out1[16], {bnn_Add_17Sx16S_17S_1_3451_out1[16], {bnn_Add_17Sx16S_17S_1_3436_out1[16], {bnn_Add_17Sx16S_17S_1_3418_out1[16], {bnn_Add_17Sx16S_17S_1_3400_out1[16], {bnn_Add_17Sx16S_17S_1_3384_out1[16], {bnn_Add_17Sx16S_17S_1_3369_out1[16], {bnn_Add_17Sx16S_17S_1_3355_out1[16], {bnn_Add_17Sx16S_17S_1_3342_out1[16]
                            , {bnn_Add_17Sx16S_17S_1_3329_out1[16], {bnn_Add_17Sx16S_17S_1_3233_out1[16], {bnn_Add_17Sx16S_17S_1_3220_out1[16], {bnn_Add_17Sx16S_17S_1_3207_out1[16], {bnn_Add_17Sx16S_17S_1_3192_out1[16], {bnn_Add_17Sx16S_17S_1_3174_out1[16], {bnn_Add_17Sx16S_17S_1_3155_out1[16], {bnn_Add_17Sx16S_17S_1_3137_out1[16], {bnn_Add_17Sx16S_17S_1_3097_out1[16], {bnn_Add_17Sx16S_17S_1_3296_out1[16], {bnn_Add_17Sx16S_17S_1_3262_out1[16], {bnn_Add_17Sx16S_17S_1_3247_out1[16]
                            , {bnn_Add_17Sx16S_17S_1_3278_out1[16], {bnn_Add_17Sx16S_17S_1_3314_out1[16], {bnn_Add_17Sx16S_17S_1_3118_out1[16], {bnn_Add_17Sx16S_17S_1_3162_out1[16], bnn_Add_17Sx16S_17S_1_2389_out1[16]}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}};
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_69bx2i
         // resource: regr_69b
         always @(posedge clk)
          begin :drive_xcelresp_data
            if (stall0) begin
            end
            else begin
               if (en_1) begin
                  case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                     7'd001: begin
                        xcelresp_data <= {bnn_N_MuxB_160_2_0_4_37_out1[139:135], 64'd00000000000000000000};
                     end
                     
                     default: begin
                        xcelresp_data <= {bnn_N_MuxB_160_2_0_4_37_out1[139:135], bnn_N_MuxB_64_10_5_4_74_out1};
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelreq_m_busy_req_0
            if (reset == 1'b1) begin
               xcelreq_m_busy_req_0 <= 1'd1;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state) 

                     5'd19: begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (en_0) begin
                                 if (drain3) begin
                                 end
                                 else begin
                                    xcelreq_m_busy_req_0 <= 1'd0;
                                 end
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (en_0) begin
                                       if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                          xcelreq_m_busy_req_0 <= 1'd1;
                                       end
                                       else begin
                                          xcelreq_m_busy_req_0 <= 1'd0;
                                       end
                                    end
                                    else begin
                                       xcelreq_m_busy_req_0 <= 1'd1;
                                    end
                                 end
                                 
                                 default: begin
                                    if (en_0) begin
                                       if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                          xcelreq_m_busy_req_0 <= 1'd1;
                                       end
                                       else begin
                                          xcelreq_m_busy_req_0 <= 1'd0;
                                       end
                                    end
                                    else begin
                                       xcelreq_m_busy_req_0 <= 1'd1;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (en_0) begin
                              if (drain3) begin
                              end
                              else begin
                                 xcelreq_m_busy_req_0 <= 1'd0;
                              end
                           end
                        end
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         always @(stall0 or en_0 or gs_ctrl4)
          begin :drive_xcelreq_m_stalling
            if (stall0) begin
               xcelreq_m_stalling = 1'd1;
            end
            else begin
               if (gs_ctrl4) begin
                  if (en_0) begin
                     xcelreq_m_stalling = 1'd0;
                  end
                  else begin
                     xcelreq_m_stalling = 1'd1;
                  end
               end
               else begin
                  xcelreq_m_stalling = 1'd0;
               end
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelresp_m_req_m_trig_req
            if (reset == 1'b1) begin
               xcelresp_m_req_m_trig_req <= 1'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state) 

                     5'd19: begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                           end
                           else begin
                              xcelresp_m_req_m_trig_req <= bnn_Not_1U_1U_4_19_out1;
                           end
                        end
                     end
                     
                  endcase

               end
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memreq_m_req_m_trig_req
            if (reset == 1'b1) begin
               memreq_m_req_m_trig_req <= 1'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state) 

                     5'd01, 5'd02: begin
                        if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                     end
                     
                     5'd04: begin
                        memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                     end
                     
                     5'd11: begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                           end
                        end
                     end
                     
                     5'd12: begin
                        if (bnn_LessThan_10Ux32U_1U_4_4104_out1) begin
                           if (3'd0 == bnn_N_Mux_3_2_6_4_4105_out1) begin
                              memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                           end
                        end
                        else begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                     end
                     
                     5'd14: begin
                        if (32'd0000000000 == s_reg_1000) begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                     end
                     
                     5'd15: begin
                        if (!cycle3_state && !s_reg_1044_stage2) begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                        else begin
                           if (cycle1_state0) begin
                           end
                           else begin
                              memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                           end
                        end
                     end
                     
                     5'd16: begin
                        if (!cycle2_state1 && !s_reg_907) begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                        else begin
                           if (cycle1_state1) begin
                              if (drain) begin
                              end
                              else begin
                                 memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                              end
                           end
                           else begin
                              if (bnn_Equal_1Ux1U_1U_1_1_4_out1) begin
                              end
                              else begin
                                 memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                              end
                           end
                        end
                     end
                     
                     5'd18: begin
                        if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                           if (s_reg_907) begin
                           end
                           else begin
                              memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                           end
                        end
                        else begin
                           memreq_m_req_m_trig_req <= bnn_Not_1U_1U_4_23_out1;
                        end
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memresp_m_busy_req_0
            if (reset == 1'b1) begin
               memresp_m_busy_req_0 <= 1'd1;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state) 

                     5'd07, 5'd13, 5'd17: begin
                        memresp_m_busy_req_0 <= 1'd0;
                     end
                     
                     5'd08, 5'd14, 5'd18: begin
                        memresp_m_busy_req_0 <= 1'd1;
                     end
                     
                     5'd11: begin
                        if (cycle1_state) begin
                           if (cycle2_state) begin
                           end
                           else begin
                              memresp_m_busy_req_0 <= 1'd1;
                           end
                        end
                        else begin
                           memresp_m_busy_req_0 <= 1'd0;
                        end
                     end
                     
                     5'd15: begin
                        if (cycle2_state0) begin
                           if (cycle3_state) begin
                           end
                           else begin
                              memresp_m_busy_req_0 <= 1'd1;
                           end
                        end
                        else begin
                           memresp_m_busy_req_0 <= 1'd0;
                        end
                     end
                     
                     5'd16: begin
                        if (cycle1_state1) begin
                           if (cycle2_state1) begin
                           end
                           else begin
                              memresp_m_busy_req_0 <= 1'd1;
                           end
                        end
                        else begin
                           memresp_m_busy_req_0 <= 1'd0;
                        end
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx4i
         always @(bnn_And_1Sx1U_1U_4_22_out1 or bnn_Not_1U_1U_4_31_out1 or cycle1_state or cycle2_state or cycle2_state0 or cycle3_state or cycle1_state1 or cycle2_state1 or global_state)
          begin :drive_stall0
            case (global_state) 

               5'd07, 5'd13, 5'd17: begin
                  stall0 = bnn_And_1Sx1U_1U_4_22_out1;
               end
               
               5'd08, 5'd14, 5'd18: begin
                  stall0 = bnn_Not_1U_1U_4_31_out1;
               end
               
               5'd11: begin
                  if (cycle2_state) begin
                     if (cycle1_state) begin
                        stall0 = 1'b0;
                     end
                     else begin
                        stall0 = bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
                  else begin
                     if (cycle1_state) begin
                        stall0 = bnn_Not_1U_1U_4_31_out1;
                     end
                     else begin
                        stall0 = bnn_Not_1U_1U_4_31_out1 | bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
               end
               
               5'd15: begin
                  if (cycle3_state) begin
                     if (cycle2_state0) begin
                        stall0 = 1'b0;
                     end
                     else begin
                        stall0 = bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
                  else begin
                     if (cycle2_state0) begin
                        stall0 = bnn_Not_1U_1U_4_31_out1;
                     end
                     else begin
                        stall0 = bnn_Not_1U_1U_4_31_out1 | bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
               end
               
               5'd16: begin
                  if (cycle2_state1) begin
                     if (cycle1_state1) begin
                        stall0 = 1'b0;
                     end
                     else begin
                        stall0 = bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
                  else begin
                     if (cycle1_state1) begin
                        stall0 = bnn_Not_1U_1U_4_31_out1;
                     end
                     else begin
                        stall0 = bnn_Not_1U_1U_4_31_out1 | bnn_And_1Sx1U_1U_4_22_out1;
                     end
                  end
               end
               
               default: begin
                  stall0 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(gs_ctrl690)
          begin :drive_fixed_buffer_0_if_0_wen0_wire
            if (gs_ctrl690) begin
               fixed_buffer_0_if_0_wen0_wire = 1'b1;
            end
            else begin
               fixed_buffer_0_if_0_wen0_wire = 1'b0;
            end
         end

         // resource: mux_4bx2i
         always @(s_reg_871[3:0] or gs_ctrl691)
          begin :drive_in1_waddr_wire
            if (gs_ctrl691) begin
               in1_waddr_wire = s_reg_871[3:0];
            end
            else begin
               in1_waddr_wire = 4'd00;
            end
         end

         // resource: mux_4bx4i
         always @(drain or drain1 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or s_reg_1034_stage1[3:0] or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl692)
          begin :drive_in1_raddr_wire
            case (gs_ctrl692) 

               3'd1: begin
                  in1_raddr_wire = 4'd00;
               end
               
               3'd2: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire = 4'd00;
                     end
                     else begin
                        in1_raddr_wire = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire = s_reg_871[3:0];
                  end
               end
               
               3'd3: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire = 4'd00;
                     end
                     else begin
                        in1_raddr_wire = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire = s_reg_1034_stage1[3:0];
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1059_stage1 or cycle2_state or gs_ctrl197)
          begin :drive_fixed_buffer_0_if_2_wen0_wire
            if (gs_ctrl197) begin
               if (!cycle2_state && s_reg_1059_stage1) begin
                  fixed_buffer_0_if_2_wen0_wire = 1'b1;
               end
               else begin
                  fixed_buffer_0_if_2_wen0_wire = 1'b0;
               end
            end
            else begin
               fixed_buffer_0_if_2_wen0_wire = 1'b0;
            end
         end

         assign in1_din_wire = bnn_Add_17Sx16S_17S_1_2389_out1[11:0];

         assign in2_waddr_wire = s_reg_1034_stage1[3:0];

         assign in1_din_wire_0 = bnn_Add_17Sx16S_17S_1_2390_out1[11:0];

         assign in1_din_wire_1 = bnn_Add_17Sx16S_17S_1_2417_out1[11:0];

         assign in1_din_wire_2 = bnn_Add_17Sx16S_17S_1_2444_out1[11:0];

         assign in1_din_wire_3 = bnn_Add_17Sx16S_17S_1_2471_out1[11:0];

         assign in1_din_wire_4 = bnn_Add_17Sx16S_17S_1_2498_out1[11:0];

         assign in1_din_wire_5 = bnn_Add_17Sx16S_17S_1_2525_out1[11:0];

         assign in1_din_wire_6 = bnn_Add_17Sx16S_17S_1_2552_out1[11:0];

         assign in1_din_wire_7 = bnn_Add_17Sx16S_17S_1_2579_out1[11:0];

         assign in1_din_wire_8 = bnn_Add_17Sx16S_17S_1_2606_out1[11:0];

         assign in1_din_wire_9 = bnn_Add_17Sx16S_17S_1_2633_out1[11:0];

         assign in1_din_wire_10 = bnn_Add_17Sx16S_17S_1_2660_out1[11:0];

         assign in1_din_wire_11 = bnn_Add_17Sx16S_17S_1_2687_out1[11:0];

         assign in1_din_wire_12 = bnn_Add_17Sx16S_17S_1_2714_out1[11:0];

         assign in1_din_wire_13 = bnn_Add_17Sx16S_17S_1_2741_out1[11:0];

         assign in1_din_wire_14 = bnn_Add_17Sx16S_17S_1_2769_out1[11:0];

         assign in1_din_wire_15 = bnn_Add_17Sx16S_17S_1_2797_out1[11:0];

         assign in1_din_wire_16 = bnn_Add_17Sx16S_17S_1_2824_out1[11:0];

         assign in1_din_wire_17 = bnn_Add_17Sx16S_17S_1_2851_out1[11:0];

         assign in1_din_wire_18 = bnn_Add_17Sx16S_17S_1_2878_out1[11:0];

         assign in1_din_wire_19 = bnn_Add_17Sx16S_17S_1_2905_out1[11:0];

         assign in1_din_wire_20 = bnn_Add_17Sx16S_17S_1_2932_out1[11:0];

         assign in1_din_wire_21 = bnn_Add_17Sx16S_17S_1_2957_out1[11:0];

         assign in1_din_wire_22 = bnn_Add_17Sx16S_17S_1_2981_out1[11:0];

         assign in1_din_wire_23 = bnn_Add_17Sx16S_17S_1_3005_out1[11:0];

         assign in1_din_wire_24 = bnn_Add_17Sx16S_17S_1_3030_out1[11:0];

         assign in1_din_wire_25 = bnn_Add_17Sx16S_17S_1_3057_out1[11:0];

         assign in1_din_wire_26 = bnn_Add_17Sx16S_17S_1_3083_out1[11:0];

         assign in1_din_wire_27 = bnn_Add_17Sx16S_17S_1_3107_out1[11:0];

         assign in1_din_wire_28 = bnn_Add_17Sx16S_17S_1_3128_out1[11:0];

         assign in1_din_wire_29 = bnn_Add_17Sx16S_17S_1_3146_out1[11:0];

         assign in1_din_wire_30 = bnn_Add_17Sx16S_17S_1_3162_out1[11:0];

         // resource: mux_4bx5i
         always @(drain or drain1 or s_reg_1013 or s_reg_1026 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl820)
          begin :drive_in1_raddr_wire_31
            case (gs_ctrl820) 

               3'd1: begin
                  in1_raddr_wire_31 = s_reg_1013;
               end
               
               3'd2: begin
                  in1_raddr_wire_31 = 4'd00;
               end
               
               3'd3: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire_31 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_31 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_31 = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire_31 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_31 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_31 = s_reg_871[3:0];
                  end
               end
               
               3'd5: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire_31 = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire_31 = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire_31 = s_reg_1026;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1034_stage1 or cycle2_state or gs_ctrl196)
          begin :drive_fixed_buffer_32_if_2_wen0_wire
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && s_reg_1034_stage1 != 10'd0000) begin
                     fixed_buffer_32_if_2_wen0_wire = 1'b1;
                  end
                  else begin
                     fixed_buffer_32_if_2_wen0_wire = 1'b0;
                  end
               end
               
               2'd2: begin
                  fixed_buffer_32_if_2_wen0_wire = 1'b1;
               end
               
               default: begin
                  fixed_buffer_32_if_2_wen0_wire = 1'b0;
               end
               
            endcase

         end

         assign in1_din_wire_31 = bnn_Add_17Sx16S_17S_1_3097_out1[11:0];

         // resource: mux_4bx2i
         always @(s_reg_1013 or bnn_Sub_4Ux1U_4S_4_1597_out1 or gs_ctrl105)
          begin :drive_in2_waddr_wire_31
            if (gs_ctrl105) begin
               in2_waddr_wire_31 = s_reg_1013;
            end
            else begin
               in2_waddr_wire_31 = bnn_Sub_4Ux1U_4S_4_1597_out1;
            end
         end

         assign in1_din_wire_32 = bnn_Add_17Sx16S_17S_1_3118_out1[11:0];

         assign in1_din_wire_33 = bnn_Add_17Sx16S_17S_1_3137_out1[11:0];

         assign in1_din_wire_34 = bnn_Add_17Sx16S_17S_1_3155_out1[11:0];

         assign in1_din_wire_35 = bnn_Add_17Sx16S_17S_1_3174_out1[11:0];

         assign in1_din_wire_36 = bnn_Add_17Sx16S_17S_1_3192_out1[11:0];

         assign in1_din_wire_37 = bnn_Add_17Sx16S_17S_1_3207_out1[11:0];

         assign in1_din_wire_38 = bnn_Add_17Sx16S_17S_1_3220_out1[11:0];

         assign in1_din_wire_39 = bnn_Add_17Sx16S_17S_1_3233_out1[11:0];

         assign in1_din_wire_40 = bnn_Add_17Sx16S_17S_1_3247_out1[11:0];

         assign in1_din_wire_41 = bnn_Add_17Sx16S_17S_1_3262_out1[11:0];

         assign in1_din_wire_42 = bnn_Add_17Sx16S_17S_1_3278_out1[11:0];

         assign in1_din_wire_43 = bnn_Add_17Sx16S_17S_1_3296_out1[11:0];

         assign in1_din_wire_44 = bnn_Add_17Sx16S_17S_1_3314_out1[11:0];

         assign in1_din_wire_45 = bnn_Add_17Sx16S_17S_1_3329_out1[11:0];

         assign in1_din_wire_46 = bnn_Add_17Sx16S_17S_1_3342_out1[11:0];

         assign in1_din_wire_47 = bnn_Add_17Sx16S_17S_1_3355_out1[11:0];

         assign in1_din_wire_48 = bnn_Add_17Sx16S_17S_1_3369_out1[11:0];

         // resource: mux_4bx5i
         always @(drain or drain1 or s_reg_1026 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or bnn_N_Mux_4_2_11_4_4090_out1 or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl820)
          begin :drive_in1_raddr_wire_49
            case (gs_ctrl820) 

               3'd1: begin
                  in1_raddr_wire_49 = bnn_N_Mux_4_2_11_4_4090_out1;
               end
               
               3'd2: begin
                  in1_raddr_wire_49 = 4'd00;
               end
               
               3'd3: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire_49 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_49 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_49 = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire_49 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_49 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_49 = s_reg_871[3:0];
                  end
               end
               
               3'd5: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire_49 = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire_49 = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire_49 = s_reg_1026;
               end
               
            endcase

         end

         assign in1_din_wire_49 = bnn_Add_17Sx16S_17S_1_3384_out1[11:0];

         // resource: mux_4bx2i
         always @(bnn_Sub_4Ux1U_4S_4_1597_out1 or bnn_N_Mux_4_2_11_4_4090_out1 or gs_ctrl105)
          begin :drive_in2_waddr_wire_49
            if (gs_ctrl105) begin
               in2_waddr_wire_49 = bnn_N_Mux_4_2_11_4_4090_out1;
            end
            else begin
               in2_waddr_wire_49 = bnn_Sub_4Ux1U_4S_4_1597_out1;
            end
         end

         assign in1_din_wire_50 = bnn_Add_17Sx16S_17S_1_3400_out1[11:0];

         assign in1_din_wire_51 = bnn_Add_17Sx16S_17S_1_3418_out1[11:0];

         assign in1_din_wire_52 = bnn_Add_17Sx16S_17S_1_3436_out1[11:0];

         assign in1_din_wire_53 = bnn_Add_17Sx16S_17S_1_3451_out1[11:0];

         assign in1_din_wire_54 = bnn_Add_17Sx16S_17S_1_3464_out1[11:0];

         assign in1_din_wire_55 = bnn_Add_17Sx16S_17S_1_3477_out1[11:0];

         assign in1_din_wire_56 = bnn_Add_17Sx16S_17S_1_3491_out1[11:0];

         // resource: mux_4bx5i
         always @(drain or drain1 or s_reg_1026 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or bnn_N_Mux_4_2_11_4_4098_out1 or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl820)
          begin :drive_in1_raddr_wire_57
            case (gs_ctrl820) 

               3'd1: begin
                  in1_raddr_wire_57 = bnn_N_Mux_4_2_11_4_4098_out1;
               end
               
               3'd2: begin
                  in1_raddr_wire_57 = 4'd00;
               end
               
               3'd3: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire_57 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_57 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_57 = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire_57 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_57 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_57 = s_reg_871[3:0];
                  end
               end
               
               3'd5: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire_57 = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire_57 = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire_57 = s_reg_1026;
               end
               
            endcase

         end

         assign in1_din_wire_57 = bnn_Add_17Sx16S_17S_1_3506_out1[11:0];

         // resource: mux_4bx2i
         always @(bnn_Sub_4Ux1U_4S_4_1597_out1 or bnn_N_Mux_4_2_11_4_4098_out1 or gs_ctrl105)
          begin :drive_in2_waddr_wire_57
            if (gs_ctrl105) begin
               in2_waddr_wire_57 = bnn_N_Mux_4_2_11_4_4098_out1;
            end
            else begin
               in2_waddr_wire_57 = bnn_Sub_4Ux1U_4S_4_1597_out1;
            end
         end

         // resource: mux_4bx5i
         always @(drain or drain1 or s_reg_1026 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or bnn_N_Mux_4_2_11_4_4099_out1 or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl820)
          begin :drive_in1_raddr_wire_58
            case (gs_ctrl820) 

               3'd1: begin
                  in1_raddr_wire_58 = bnn_N_Mux_4_2_11_4_4099_out1;
               end
               
               3'd2: begin
                  in1_raddr_wire_58 = 4'd00;
               end
               
               3'd3: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire_58 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_58 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_58 = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire_58 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_58 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_58 = s_reg_871[3:0];
                  end
               end
               
               3'd5: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire_58 = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire_58 = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire_58 = s_reg_1026;
               end
               
            endcase

         end

         assign in1_din_wire_58 = bnn_Add_17Sx16S_17S_1_3521_out1[11:0];

         // resource: mux_4bx2i
         always @(bnn_Sub_4Ux1U_4S_4_1597_out1 or bnn_N_Mux_4_2_11_4_4099_out1 or gs_ctrl105)
          begin :drive_in2_waddr_wire_58
            if (gs_ctrl105) begin
               in2_waddr_wire_58 = bnn_N_Mux_4_2_11_4_4099_out1;
            end
            else begin
               in2_waddr_wire_58 = bnn_Sub_4Ux1U_4S_4_1597_out1;
            end
         end

         // resource: mux_4bx5i
         always @(drain or drain1 or s_reg_1026 or s_reg_871[3:0] or s_reg_886[3:0] or s_reg_907 or bnn_Add_7Sx5S_7S_4_195_out1[6] or bnn_N_Mux_4_2_11_4_4100_out1 or s_reg_1044_stage2 or cycle3_state or cycle2_state1 or gs_ctrl820)
          begin :drive_in1_raddr_wire_59
            case (gs_ctrl820) 

               3'd1: begin
                  in1_raddr_wire_59 = bnn_N_Mux_4_2_11_4_4100_out1;
               end
               
               3'd2: begin
                  in1_raddr_wire_59 = 4'd00;
               end
               
               3'd3: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        in1_raddr_wire_59 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_59 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_59 = s_reg_871[3:0];
                  end
               end
               
               3'd4: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     if (drain) begin
                        in1_raddr_wire_59 = 4'd00;
                     end
                     else begin
                        in1_raddr_wire_59 = s_reg_871[3:0];
                     end
                  end
                  else begin
                     in1_raddr_wire_59 = s_reg_871[3:0];
                  end
               end
               
               3'd5: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     in1_raddr_wire_59 = s_reg_886[3:0];
                  end
                  else begin
                     in1_raddr_wire_59 = s_reg_871[3:0];
                  end
               end
               
               default: begin
                  in1_raddr_wire_59 = s_reg_1026;
               end
               
            endcase

         end

         assign in1_din_wire_59 = bnn_Add_17Sx16S_17S_1_3534_out1[11:0];

         // resource: mux_4bx2i
         always @(bnn_Sub_4Ux1U_4S_4_1597_out1 or bnn_N_Mux_4_2_11_4_4100_out1 or gs_ctrl105)
          begin :drive_in2_waddr_wire_59
            if (gs_ctrl105) begin
               in2_waddr_wire_59 = bnn_N_Mux_4_2_11_4_4100_out1;
            end
            else begin
               in2_waddr_wire_59 = bnn_Sub_4Ux1U_4S_4_1597_out1;
            end
         end

         assign in1_din_wire_60 = bnn_Add_17Sx16S_17S_1_3542_out1[11:0];

         assign in1_din_wire_61 = bnn_Add_17Sx16S_17S_1_3546_out1[11:0];

         assign in1_din_wire_62 = bnn_Add_17Sx16S_17S_1_3547_out1[11:0];

         // resource: mux_2bx2i
         always @(s_reg_887 or cycle2_state or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :drive_Bline_buffer_0_mi61
            if (cycle2_state) begin
               Bline_buffer_0_mi61 = s_reg_887;
            end
            else begin
               Bline_buffer_0_mi61 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_874[1:0] or bnn_N_Mux_2_2_3_1_1831_out1 or cycle2_state)
          begin :drive_Bline_buffer_1_mi61
            if (cycle2_state) begin
               Bline_buffer_1_mi61 = s_reg_874[1:0];
            end
            else begin
               Bline_buffer_1_mi61 = bnn_N_Mux_2_2_3_1_1831_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_875 or bnn_N_Mux_2_2_3_1_1846_out1 or cycle2_state)
          begin :drive_Bline_buffer_2_mi61
            if (cycle2_state) begin
               Bline_buffer_2_mi61 = s_reg_875;
            end
            else begin
               Bline_buffer_2_mi61 = bnn_N_Mux_2_2_3_1_1846_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_881 or bnn_N_Mux_2_2_3_1_1857_out1 or cycle2_state)
          begin :drive_Bline_buffer_3_mi61
            if (cycle2_state) begin
               Bline_buffer_3_mi61 = s_reg_881;
            end
            else begin
               Bline_buffer_3_mi61 = bnn_N_Mux_2_2_3_1_1857_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_888 or bnn_N_Mux_2_2_3_1_1868_out1 or cycle2_state)
          begin :drive_Bline_buffer_4_mi61
            if (cycle2_state) begin
               Bline_buffer_4_mi61 = s_reg_888;
            end
            else begin
               Bline_buffer_4_mi61 = bnn_N_Mux_2_2_3_1_1868_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_876 or bnn_N_Mux_64_2_2_1_1636_out1[32] or cycle2_state)
          begin :drive_Bline_buffer_11_mi61
            if (cycle2_state) begin
               Bline_buffer_11_mi61 = s_reg_876;
            end
            else begin
               Bline_buffer_11_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_898 or bnn_N_Mux_2_2_3_1_1879_out1 or cycle2_state)
          begin :drive_Bline_buffer_5_mi61
            if (cycle2_state) begin
               Bline_buffer_5_mi61 = s_reg_898;
            end
            else begin
               Bline_buffer_5_mi61 = bnn_N_Mux_2_2_3_1_1879_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_877 or bnn_N_Mux_64_2_2_1_1636_out1[33] or cycle2_state)
          begin :drive_Bline_buffer_12_mi61
            if (cycle2_state) begin
               Bline_buffer_12_mi61 = s_reg_877;
            end
            else begin
               Bline_buffer_12_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_909 or bnn_N_Mux_2_2_3_1_1890_out1 or cycle2_state)
          begin :drive_Bline_buffer_6_mi61
            if (cycle2_state) begin
               Bline_buffer_6_mi61 = s_reg_909;
            end
            else begin
               Bline_buffer_6_mi61 = bnn_N_Mux_2_2_3_1_1890_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_882 or bnn_N_Mux_64_2_2_1_1636_out1[34] or cycle2_state)
          begin :drive_Bline_buffer_13_mi61
            if (cycle2_state) begin
               Bline_buffer_13_mi61 = s_reg_882;
            end
            else begin
               Bline_buffer_13_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[34], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_883 or cycle2_state or bnn_N_Mux_3_2_6_4_2178_out1_slice)
          begin :drive_Bline_buffer_20_mi61
            if (cycle2_state) begin
               Bline_buffer_20_mi61 = s_reg_883;
            end
            else begin
               Bline_buffer_20_mi61 = bnn_N_Mux_3_2_6_4_2178_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_917 or bnn_N_Mux_2_2_3_1_1901_out1 or cycle2_state)
          begin :drive_Bline_buffer_7_mi61
            if (cycle2_state) begin
               Bline_buffer_7_mi61 = s_reg_917;
            end
            else begin
               Bline_buffer_7_mi61 = bnn_N_Mux_2_2_3_1_1901_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_889 or bnn_N_Mux_64_2_2_1_1636_out1[35] or cycle2_state)
          begin :drive_Bline_buffer_14_mi61
            if (cycle2_state) begin
               Bline_buffer_14_mi61 = s_reg_889;
            end
            else begin
               Bline_buffer_14_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_925 or bnn_N_Mux_2_2_3_1_1912_out1 or cycle2_state)
          begin :drive_Bline_buffer_8_mi61
            if (cycle2_state) begin
               Bline_buffer_8_mi61 = s_reg_925;
            end
            else begin
               Bline_buffer_8_mi61 = bnn_N_Mux_2_2_3_1_1912_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_899 or bnn_N_Mux_64_2_2_1_1636_out1[36] or cycle2_state)
          begin :drive_Bline_buffer_15_mi61
            if (cycle2_state) begin
               Bline_buffer_15_mi61 = s_reg_899;
            end
            else begin
               Bline_buffer_15_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_933 or bnn_N_Mux_2_2_3_1_2164_out1 or cycle2_state)
          begin :drive_Bline_buffer_9_mi61
            if (cycle2_state) begin
               Bline_buffer_9_mi61 = s_reg_933;
            end
            else begin
               Bline_buffer_9_mi61 = bnn_N_Mux_2_2_3_1_2164_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_910 or bnn_N_Mux_64_2_2_1_1636_out1[37] or cycle2_state)
          begin :drive_Bline_buffer_16_mi61
            if (cycle2_state) begin
               Bline_buffer_16_mi61 = s_reg_910;
            end
            else begin
               Bline_buffer_16_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[37], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_891 or bnn_N_Mux_2_2_3_1_2176_out1 or cycle2_state)
          begin :drive_Bline_buffer_30_mi61
            if (cycle2_state) begin
               Bline_buffer_30_mi61 = s_reg_891;
            end
            else begin
               Bline_buffer_30_mi61 = bnn_N_Mux_2_2_3_1_2176_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_879 or bnn_N_Mux_2_2_3_1_1933_out1 or cycle2_state)
          begin :drive_Bline_buffer_31_mi61
            if (cycle2_state) begin
               Bline_buffer_31_mi61 = s_reg_879;
            end
            else begin
               Bline_buffer_31_mi61 = bnn_N_Mux_2_2_3_1_1933_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_918 or bnn_N_Mux_64_2_2_1_1636_out1[38] or cycle2_state)
          begin :drive_Bline_buffer_17_mi61
            if (cycle2_state) begin
               Bline_buffer_17_mi61 = s_reg_918;
            end
            else begin
               Bline_buffer_17_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[38], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_880 or bnn_N_Mux_2_2_3_1_1944_out1 or cycle2_state)
          begin :drive_Bline_buffer_32_mi61
            if (cycle2_state) begin
               Bline_buffer_32_mi61 = s_reg_880;
            end
            else begin
               Bline_buffer_32_mi61 = bnn_N_Mux_2_2_3_1_1944_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_926 or bnn_N_Mux_64_2_2_1_1636_out1[39] or cycle2_state)
          begin :drive_Bline_buffer_18_mi61
            if (cycle2_state) begin
               Bline_buffer_18_mi61 = s_reg_926;
            end
            else begin
               Bline_buffer_18_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[39], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_885 or bnn_N_Mux_2_2_3_1_1955_out1 or cycle2_state)
          begin :drive_Bline_buffer_33_mi61
            if (cycle2_state) begin
               Bline_buffer_33_mi61 = s_reg_885;
            end
            else begin
               Bline_buffer_33_mi61 = bnn_N_Mux_2_2_3_1_1955_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_902 or cycle2_state or bnn_N_Mux_3_2_6_4_1638_out1_slice)
          begin :drive_Bline_buffer_40_mi61
            if (cycle2_state) begin
               Bline_buffer_40_mi61 = s_reg_902;
            end
            else begin
               Bline_buffer_40_mi61 = bnn_N_Mux_3_2_6_4_1638_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_934 or cycle2_state or bnn_N_Mux_3_2_6_4_1637_out1_slice)
          begin :drive_Bline_buffer_19_mi61
            if (cycle2_state) begin
               Bline_buffer_19_mi61 = s_reg_934;
            end
            else begin
               Bline_buffer_19_mi61 = bnn_N_Mux_3_2_6_4_1637_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_892 or bnn_N_Mux_2_2_3_1_1966_out1 or cycle2_state)
          begin :drive_Bline_buffer_34_mi61
            if (cycle2_state) begin
               Bline_buffer_34_mi61 = s_reg_892;
            end
            else begin
               Bline_buffer_34_mi61 = bnn_N_Mux_2_2_3_1_1966_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_893 or bnn_N_Mux_64_2_2_1_1636_out1[40] or cycle2_state)
          begin :drive_Bline_buffer_41_mi61
            if (cycle2_state) begin
               Bline_buffer_41_mi61 = s_reg_893;
            end
            else begin
               Bline_buffer_41_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_901 or bnn_N_Mux_2_2_3_1_1977_out1 or cycle2_state)
          begin :drive_Bline_buffer_35_mi61
            if (cycle2_state) begin
               Bline_buffer_35_mi61 = s_reg_901;
            end
            else begin
               Bline_buffer_35_mi61 = bnn_N_Mux_2_2_3_1_1977_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_903 or bnn_N_Mux_64_2_2_1_1636_out1[41] or cycle2_state)
          begin :drive_Bline_buffer_42_mi61
            if (cycle2_state) begin
               Bline_buffer_42_mi61 = s_reg_903;
            end
            else begin
               Bline_buffer_42_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_912 or bnn_N_Mux_2_2_3_1_1988_out1 or cycle2_state)
          begin :drive_Bline_buffer_36_mi61
            if (cycle2_state) begin
               Bline_buffer_36_mi61 = s_reg_912;
            end
            else begin
               Bline_buffer_36_mi61 = bnn_N_Mux_2_2_3_1_1988_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_913 or bnn_N_Mux_64_2_2_1_1636_out1[42] or cycle2_state)
          begin :drive_Bline_buffer_43_mi61
            if (cycle2_state) begin
               Bline_buffer_43_mi61 = s_reg_913;
            end
            else begin
               Bline_buffer_43_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[42], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_920 or bnn_N_Mux_2_2_3_1_1999_out1 or cycle2_state)
          begin :drive_Bline_buffer_37_mi61
            if (cycle2_state) begin
               Bline_buffer_37_mi61 = s_reg_920;
            end
            else begin
               Bline_buffer_37_mi61 = bnn_N_Mux_2_2_3_1_1999_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_921 or bnn_N_Mux_64_2_2_1_1636_out1[43] or cycle2_state)
          begin :drive_Bline_buffer_44_mi61
            if (cycle2_state) begin
               Bline_buffer_44_mi61 = s_reg_921;
            end
            else begin
               Bline_buffer_44_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[43], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_928 or bnn_N_Mux_2_2_3_1_2010_out1 or cycle2_state)
          begin :drive_Bline_buffer_38_mi61
            if (cycle2_state) begin
               Bline_buffer_38_mi61 = s_reg_928;
            end
            else begin
               Bline_buffer_38_mi61 = bnn_N_Mux_2_2_3_1_2010_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_929 or bnn_N_Mux_64_2_2_1_1636_out1[44] or cycle2_state)
          begin :drive_Bline_buffer_45_mi61
            if (cycle2_state) begin
               Bline_buffer_45_mi61 = s_reg_929;
            end
            else begin
               Bline_buffer_45_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[44], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_935 or bnn_N_Mux_2_2_3_1_2190_out1 or cycle2_state)
          begin :drive_Bline_buffer_39_mi61
            if (cycle2_state) begin
               Bline_buffer_39_mi61 = s_reg_935;
            end
            else begin
               Bline_buffer_39_mi61 = bnn_N_Mux_2_2_3_1_2190_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_936 or bnn_N_Mux_64_2_2_1_1636_out1[45] or cycle2_state)
          begin :drive_Bline_buffer_46_mi61
            if (cycle2_state) begin
               Bline_buffer_46_mi61 = s_reg_936;
            end
            else begin
               Bline_buffer_46_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_905 or bnn_N_Mux_2_2_3_1_2208_out1 or cycle2_state)
          begin :drive_Bline_buffer_60_mi61
            if (cycle2_state) begin
               Bline_buffer_60_mi61 = s_reg_905;
            end
            else begin
               Bline_buffer_60_mi61 = bnn_N_Mux_2_2_3_1_2208_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_896 or bnn_N_Mux_2_2_3_1_2021_out1 or cycle2_state)
          begin :drive_Bline_buffer_61_mi61
            if (cycle2_state) begin
               Bline_buffer_61_mi61 = s_reg_896;
            end
            else begin
               Bline_buffer_61_mi61 = bnn_N_Mux_2_2_3_1_2021_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_940 or bnn_N_Mux_64_2_2_1_1636_out1[46] or cycle2_state)
          begin :drive_Bline_buffer_47_mi61
            if (cycle2_state) begin
               Bline_buffer_47_mi61 = s_reg_940;
            end
            else begin
               Bline_buffer_47_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_906 or bnn_N_Mux_2_2_3_1_2038_out1 or cycle2_state)
          begin :drive_Bline_buffer_62_mi61
            if (cycle2_state) begin
               Bline_buffer_62_mi61 = s_reg_906;
            end
            else begin
               Bline_buffer_62_mi61 = bnn_N_Mux_2_2_3_1_2038_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_945 or bnn_N_Mux_64_2_2_1_1636_out1[47] or cycle2_state)
          begin :drive_Bline_buffer_48_mi61
            if (cycle2_state) begin
               Bline_buffer_48_mi61 = s_reg_945;
            end
            else begin
               Bline_buffer_48_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[47], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_915 or bnn_N_Mux_2_2_3_1_2055_out1 or cycle2_state)
          begin :drive_Bline_buffer_63_mi61
            if (cycle2_state) begin
               Bline_buffer_63_mi61 = s_reg_915;
            end
            else begin
               Bline_buffer_63_mi61 = bnn_N_Mux_2_2_3_1_2055_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_948 or cycle2_state or bnn_N_Mux_3_2_6_4_1640_out1_slice)
          begin :drive_Bline_buffer_70_mi61
            if (cycle2_state) begin
               Bline_buffer_70_mi61 = s_reg_948;
            end
            else begin
               Bline_buffer_70_mi61 = bnn_N_Mux_3_2_6_4_1640_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_952 or cycle2_state or bnn_N_Mux_3_2_6_1_1639_out1_slice)
          begin :drive_Bline_buffer_49_mi61
            if (cycle2_state) begin
               Bline_buffer_49_mi61 = s_reg_952;
            end
            else begin
               Bline_buffer_49_mi61 = bnn_N_Mux_3_2_6_1_1639_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_923 or bnn_N_Mux_2_2_3_1_2072_out1 or cycle2_state)
          begin :drive_Bline_buffer_64_mi61
            if (cycle2_state) begin
               Bline_buffer_64_mi61 = s_reg_923;
            end
            else begin
               Bline_buffer_64_mi61 = bnn_N_Mux_2_2_3_1_2072_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_954 or bnn_N_Mux_64_2_2_1_1636_out1[48] or cycle2_state)
          begin :drive_Bline_buffer_71_mi61
            if (cycle2_state) begin
               Bline_buffer_71_mi61 = s_reg_954;
            end
            else begin
               Bline_buffer_71_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[48], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_931 or bnn_N_Mux_2_2_3_1_2089_out1 or cycle2_state)
          begin :drive_Bline_buffer_65_mi61
            if (cycle2_state) begin
               Bline_buffer_65_mi61 = s_reg_931;
            end
            else begin
               Bline_buffer_65_mi61 = bnn_N_Mux_2_2_3_1_2089_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_958 or bnn_N_Mux_64_2_2_1_1636_out1[49] or cycle2_state)
          begin :drive_Bline_buffer_72_mi61
            if (cycle2_state) begin
               Bline_buffer_72_mi61 = s_reg_958;
            end
            else begin
               Bline_buffer_72_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[49], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_938 or bnn_N_Mux_2_2_3_1_2106_out1 or cycle2_state)
          begin :drive_Bline_buffer_66_mi61
            if (cycle2_state) begin
               Bline_buffer_66_mi61 = s_reg_938;
            end
            else begin
               Bline_buffer_66_mi61 = bnn_N_Mux_2_2_3_1_2106_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_961 or bnn_N_Mux_64_2_2_1_1636_out1[50] or cycle2_state)
          begin :drive_Bline_buffer_73_mi61
            if (cycle2_state) begin
               Bline_buffer_73_mi61 = s_reg_961;
            end
            else begin
               Bline_buffer_73_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[50], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_942 or bnn_N_Mux_2_2_3_1_2123_out1 or cycle2_state)
          begin :drive_Bline_buffer_67_mi61
            if (cycle2_state) begin
               Bline_buffer_67_mi61 = s_reg_942;
            end
            else begin
               Bline_buffer_67_mi61 = bnn_N_Mux_2_2_3_1_2123_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_964 or bnn_N_Mux_64_2_2_1_1636_out1[51] or cycle2_state)
          begin :drive_Bline_buffer_74_mi61
            if (cycle2_state) begin
               Bline_buffer_74_mi61 = s_reg_964;
            end
            else begin
               Bline_buffer_74_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[51], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_947 or bnn_N_Mux_2_2_3_1_2140_out1 or cycle2_state)
          begin :drive_Bline_buffer_68_mi61
            if (cycle2_state) begin
               Bline_buffer_68_mi61 = s_reg_947;
            end
            else begin
               Bline_buffer_68_mi61 = bnn_N_Mux_2_2_3_1_2140_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_967 or bnn_N_Mux_64_2_2_1_1636_out1[52] or cycle2_state)
          begin :drive_Bline_buffer_75_mi61
            if (cycle2_state) begin
               Bline_buffer_75_mi61 = s_reg_967;
            end
            else begin
               Bline_buffer_75_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[52], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_953 or bnn_N_Mux_2_2_3_1_2196_out1 or cycle2_state)
          begin :drive_Bline_buffer_69_mi61
            if (cycle2_state) begin
               Bline_buffer_69_mi61 = s_reg_953;
            end
            else begin
               Bline_buffer_69_mi61 = bnn_N_Mux_2_2_3_1_2196_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_970 or bnn_N_Mux_64_2_2_1_1636_out1[53] or cycle2_state)
          begin :drive_Bline_buffer_76_mi61
            if (cycle2_state) begin
               Bline_buffer_76_mi61 = s_reg_970;
            end
            else begin
               Bline_buffer_76_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[53], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_950 or bnn_N_Mux_2_2_3_1_2214_out1 or cycle2_state)
          begin :drive_Bline_buffer_90_mi61
            if (cycle2_state) begin
               Bline_buffer_90_mi61 = s_reg_950;
            end
            else begin
               Bline_buffer_90_mi61 = bnn_N_Mux_2_2_3_1_2214_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_956 or bnn_N_Mux_2_2_3_1_2027_out1 or cycle2_state)
          begin :drive_Bline_buffer_91_mi61
            if (cycle2_state) begin
               Bline_buffer_91_mi61 = s_reg_956;
            end
            else begin
               Bline_buffer_91_mi61 = bnn_N_Mux_2_2_3_1_2027_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_973 or bnn_N_Mux_64_2_2_1_1636_out1[54] or cycle2_state)
          begin :drive_Bline_buffer_77_mi61
            if (cycle2_state) begin
               Bline_buffer_77_mi61 = s_reg_973;
            end
            else begin
               Bline_buffer_77_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[54], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_960 or bnn_N_Mux_2_2_3_1_2044_out1 or cycle2_state)
          begin :drive_Bline_buffer_92_mi61
            if (cycle2_state) begin
               Bline_buffer_92_mi61 = s_reg_960;
            end
            else begin
               Bline_buffer_92_mi61 = bnn_N_Mux_2_2_3_1_2044_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_978 or bnn_N_Mux_64_2_2_1_1636_out1[55] or cycle2_state)
          begin :drive_Bline_buffer_78_mi61
            if (cycle2_state) begin
               Bline_buffer_78_mi61 = s_reg_978;
            end
            else begin
               Bline_buffer_78_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[55], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_963 or bnn_N_Mux_2_2_3_1_2061_out1 or cycle2_state)
          begin :drive_Bline_buffer_93_mi61
            if (cycle2_state) begin
               Bline_buffer_93_mi61 = s_reg_963;
            end
            else begin
               Bline_buffer_93_mi61 = bnn_N_Mux_2_2_3_1_2061_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_981 or cycle2_state or bnn_N_Mux_3_2_6_1_1642_out1_slice)
          begin :drive_Bline_buffer_100_mi61
            if (cycle2_state) begin
               Bline_buffer_100_mi61 = s_reg_981;
            end
            else begin
               Bline_buffer_100_mi61 = bnn_N_Mux_3_2_6_1_1642_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_983 or cycle2_state or bnn_N_Mux_3_2_6_1_1641_out1_slice)
          begin :drive_Bline_buffer_79_mi61
            if (cycle2_state) begin
               Bline_buffer_79_mi61 = s_reg_983;
            end
            else begin
               Bline_buffer_79_mi61 = bnn_N_Mux_3_2_6_1_1641_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_966 or bnn_N_Mux_2_2_3_1_2078_out1 or cycle2_state)
          begin :drive_Bline_buffer_94_mi61
            if (cycle2_state) begin
               Bline_buffer_94_mi61 = s_reg_966;
            end
            else begin
               Bline_buffer_94_mi61 = bnn_N_Mux_2_2_3_1_2078_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_985 or bnn_N_Mux_64_2_2_1_1636_out1[56] or cycle2_state)
          begin :drive_Bline_buffer_101_mi61
            if (cycle2_state) begin
               Bline_buffer_101_mi61 = s_reg_985;
            end
            else begin
               Bline_buffer_101_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[56], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_969 or bnn_N_Mux_2_2_3_1_2095_out1 or cycle2_state)
          begin :drive_Bline_buffer_95_mi61
            if (cycle2_state) begin
               Bline_buffer_95_mi61 = s_reg_969;
            end
            else begin
               Bline_buffer_95_mi61 = bnn_N_Mux_2_2_3_1_2095_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_987 or bnn_N_Mux_64_2_2_1_1636_out1[57] or cycle2_state)
          begin :drive_Bline_buffer_102_mi61
            if (cycle2_state) begin
               Bline_buffer_102_mi61 = s_reg_987;
            end
            else begin
               Bline_buffer_102_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[57], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_972 or bnn_N_Mux_2_2_3_1_2112_out1 or cycle2_state)
          begin :drive_Bline_buffer_96_mi61
            if (cycle2_state) begin
               Bline_buffer_96_mi61 = s_reg_972;
            end
            else begin
               Bline_buffer_96_mi61 = bnn_N_Mux_2_2_3_1_2112_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_989 or bnn_N_Mux_64_2_2_1_1636_out1[58] or cycle2_state)
          begin :drive_Bline_buffer_103_mi61
            if (cycle2_state) begin
               Bline_buffer_103_mi61 = s_reg_989;
            end
            else begin
               Bline_buffer_103_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[58], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_975 or bnn_N_Mux_2_2_3_1_2129_out1 or cycle2_state)
          begin :drive_Bline_buffer_97_mi61
            if (cycle2_state) begin
               Bline_buffer_97_mi61 = s_reg_975;
            end
            else begin
               Bline_buffer_97_mi61 = bnn_N_Mux_2_2_3_1_2129_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_991 or bnn_N_Mux_64_2_2_1_1636_out1[59] or cycle2_state)
          begin :drive_Bline_buffer_104_mi61
            if (cycle2_state) begin
               Bline_buffer_104_mi61 = s_reg_991;
            end
            else begin
               Bline_buffer_104_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[59], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_980 or bnn_N_Mux_2_2_3_4_2146_out1 or cycle2_state)
          begin :drive_Bline_buffer_98_mi61
            if (cycle2_state) begin
               Bline_buffer_98_mi61 = s_reg_980;
            end
            else begin
               Bline_buffer_98_mi61 = bnn_N_Mux_2_2_3_4_2146_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_993 or bnn_N_Mux_64_2_2_1_1636_out1[60] or cycle2_state)
          begin :drive_Bline_buffer_105_mi61
            if (cycle2_state) begin
               Bline_buffer_105_mi61 = s_reg_993;
            end
            else begin
               Bline_buffer_105_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[60], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_995 or bnn_N_Mux_64_2_2_1_1636_out1[61] or cycle2_state)
          begin :drive_Bline_buffer_106_mi61
            if (cycle2_state) begin
               Bline_buffer_106_mi61 = s_reg_995;
            end
            else begin
               Bline_buffer_106_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[61], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_984 or cycle2_state or bnn_N_Mux_3_2_6_4_1833_out1_slice)
          begin :drive_Bline_buffer_99_mi61
            if (cycle2_state) begin
               Bline_buffer_99_mi61 = s_reg_984;
            end
            else begin
               Bline_buffer_99_mi61 = bnn_N_Mux_3_2_6_4_1833_out1_slice;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_997 or bnn_N_Mux_64_2_2_1_1636_out1[62] or cycle2_state)
          begin :drive_Bline_buffer_107_mi61
            if (cycle2_state) begin
               Bline_buffer_107_mi61 = s_reg_997;
            end
            else begin
               Bline_buffer_107_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[62], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_999 or bnn_N_Mux_64_2_2_1_1636_out1[63] or cycle2_state)
          begin :drive_Bline_buffer_108_mi61
            if (cycle2_state) begin
               Bline_buffer_108_mi61 = s_reg_999;
            end
            else begin
               Bline_buffer_108_mi61 = {bnn_N_Mux_64_2_2_1_1636_out1[63], 1'b1};
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_977 or cycle2_state or bnn_N_Mux_3_2_6_4_1835_out1_slice)
          begin :drive_Bline_buffer_119_mi61
            if (cycle2_state) begin
               Bline_buffer_119_mi61 = s_reg_977;
            end
            else begin
               Bline_buffer_119_mi61 = bnn_N_Mux_3_2_6_4_1835_out1_slice;
            end
         end

         // resource: mux_64bx2i
         always @(bnn_N_Mux_64_2_2_1_5202_out1 or cycle1_state0)
          begin :drive_Boutword_i0_mi87
            if (cycle1_state0) begin
               Boutword_i0_mi87 = 64'd18446744073709551615;
            end
            else begin
               Boutword_i0_mi87 = bnn_N_Mux_64_2_2_1_5202_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_872 or bnn_N_Mux_2_2_3_4_62_out1 or cycle1_state2)
          begin :drive_short_width_mode_mi9
            if (cycle1_state2) begin
               short_width_mode_mi9 = s_reg_872;
            end
            else begin
               short_width_mode_mi9 = bnn_N_Mux_2_2_3_4_62_out1;
            end
         end

         // resource: mux_64bx2i
         always @(s_reg_897 or bnn_N_Mux_64_2_2_4_63_out1 or cycle1_state2)
          begin :drive_short_n_inputs_mi9
            if (cycle1_state2) begin
               short_n_inputs_mi9 = s_reg_897;
            end
            else begin
               short_n_inputs_mi9 = bnn_N_Mux_64_2_2_4_63_out1;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_870 or bnn_And_1Sx1U_1U_4_67_out1 or cycle1_state2)
          begin :drive_short_popped_go_0_u0_mi9
            if (cycle1_state2) begin
               short_popped_go_0_u0_mi9 = s_reg_870;
            end
            else begin
               short_popped_go_0_u0_mi9 = bnn_And_1Sx1U_1U_4_67_out1;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_907 or bnn_N_Muxb_1_2_18_4_68_out1 or cycle1_state2)
          begin :drive_short_do_max_pool_mi9
            if (cycle1_state2) begin
               short_do_max_pool_mi9 = s_reg_907;
            end
            else begin
               short_do_max_pool_mi9 = bnn_N_Muxb_1_2_18_4_68_out1;
            end
         end

         // resource: mux_32bx2i
         always @(s_reg_1017 or bnn_N_Mux_32_2_1_4_69_out1 or cycle1_state2)
          begin :drive_short_addr_w_mi9
            if (cycle1_state2) begin
               short_addr_w_mi9 = s_reg_1017;
            end
            else begin
               short_addr_w_mi9 = bnn_N_Mux_32_2_1_4_69_out1;
            end
         end

         // resource: mux_32bx2i
         always @(s_reg_1003 or bnn_N_Mux_32_2_1_4_70_out1 or cycle1_state2)
          begin :drive_short_addr_kh_mi9
            if (cycle1_state2) begin
               short_addr_kh_mi9 = s_reg_1003;
            end
            else begin
               short_addr_kh_mi9 = bnn_N_Mux_32_2_1_4_70_out1;
            end
         end

         // resource: mux_32bx2i
         always @(s_reg_1002 or bnn_N_Mux_32_2_1_4_71_out1 or cycle1_state2)
          begin :drive_short_addr_in_fmap_mi9
            if (cycle1_state2) begin
               short_addr_in_fmap_mi9 = s_reg_1002;
            end
            else begin
               short_addr_in_fmap_mi9 = bnn_N_Mux_32_2_1_4_71_out1;
            end
         end

         // resource: mux_32bx2i
         always @(s_reg_1001 or bnn_N_Mux_32_2_1_4_72_out1 or cycle1_state2)
          begin :drive_short_addr_out_fmap_mi9
            if (cycle1_state2) begin
               short_addr_out_fmap_mi9 = s_reg_1001;
            end
            else begin
               short_addr_out_fmap_mi9 = bnn_N_Mux_32_2_1_4_72_out1;
            end
         end

         // resource: mux_32bx2i
         always @(s_reg_1000 or bnn_N_Mux_32_2_1_4_73_out1 or cycle1_state2)
          begin :drive_short_addr_conv_out_mi9
            if (cycle1_state2) begin
               short_addr_conv_out_mi9 = s_reg_1000;
            end
            else begin
               short_addr_conv_out_mi9 = bnn_N_Mux_32_2_1_4_73_out1;
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_drain
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (!s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        drain <= 1'd0;
                     end
                  end
                  
                  5'd16: begin
                     if (cycle1_state1) begin
                     end
                     else begin
                        drain <= bnn_Equal_1Ux1U_1U_1_1_4_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_drain1
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        drain1 <= 1'd0;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                     end
                     else begin
                        drain1 <= bnn_Equal_1Ux1U_1U_1_1_3_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_drain2
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        drain2 <= 1'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        drain2 <= bnn_Equal_1Ux1U_1U_1_1_2_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_drain3
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     drain3 <= 1'd0;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        drain3 <= 1'd0;
                     end
                  end
                  
                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                              7'd001: begin
                                 drain3 <= bnn_Equal_1Ux1U_1U_1_1_1_out1;
                              end
                              
                              default: begin
                                 drain3 <= bnn_Equal_1Ux1U_1U_1_1_out1;
                              end
                              
                           endcase

                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_32bx4i
         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1000
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_1000 <= 32'd0000000000;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_1000 <= s_reg_1011;
                     end
                  end
                  
                  5'd19: begin
                     if (en_2) begin
                        case (cycle2_state2) 

                           2'd0, 2'd1: begin
                              if (s_reg_870_stage10) begin
                                 if (en_0) begin
                                    if (en_1) begin
                                       if (cycle1_state2) begin
                                          if (drain3) begin
                                          end
                                          else begin
                                             s_reg_1000 <= short_addr_conv_out_mi9;
                                          end
                                       end
                                       else begin
                                          case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                             7'd001: begin
                                                if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                                end
                                                else begin
                                                   s_reg_1000 <= short_addr_conv_out_mi9;
                                                end
                                             end
                                             
                                             default: begin
                                                if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                                end
                                                else begin
                                                   s_reg_1000 <= short_addr_conv_out_mi9;
                                                end
                                             end
                                             
                                          endcase

                                       end
                                    end
                                    else begin
                                       if (drain3) begin
                                       end
                                       else begin
                                          s_reg_1000 <= short_addr_conv_out_mi9;
                                       end
                                    end
                                 end
                              end
                              else begin
                                 if (en_0) begin
                                    if (en_1) begin
                                       if (cycle1_state2) begin
                                          if (drain3) begin
                                             /* state15 */
                                             s_reg_1000 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                                          end
                                          else begin
                                             s_reg_1000 <= short_addr_conv_out_mi9;
                                          end
                                       end
                                       else begin
                                          case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                             7'd001: begin
                                                if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                                   /* state15 */
                                                   s_reg_1000 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                                                end
                                                else begin
                                                   s_reg_1000 <= short_addr_conv_out_mi9;
                                                end
                                             end
                                             
                                             default: begin
                                                if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                                   /* state15 */
                                                   s_reg_1000 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                                                end
                                                else begin
                                                   s_reg_1000 <= short_addr_conv_out_mi9;
                                                end
                                             end
                                             
                                          endcase

                                       end
                                    end
                                    else begin
                                       if (drain3) begin
                                          /* state15 */
                                          s_reg_1000 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                                       end
                                       else begin
                                          s_reg_1000 <= short_addr_conv_out_mi9;
                                       end
                                    end
                                 end
                                 else begin
                                    /* state15 */
                                    s_reg_1000 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                                 end
                              end
                           end
                           
                           default: begin
                              if (en_0) begin
                                 if (en_1) begin
                                    if (cycle1_state2) begin
                                       if (drain3) begin
                                       end
                                       else begin
                                          s_reg_1000 <= short_addr_conv_out_mi9;
                                       end
                                    end
                                    else begin
                                       case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                          7'd001: begin
                                             if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                             end
                                             else begin
                                                s_reg_1000 <= short_addr_conv_out_mi9;
                                             end
                                          end
                                          
                                          default: begin
                                             if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                             end
                                             else begin
                                                s_reg_1000 <= short_addr_conv_out_mi9;
                                             end
                                          end
                                          
                                       endcase

                                    end
                                 end
                                 else begin
                                    if (drain3) begin
                                    end
                                    else begin
                                       s_reg_1000 <= short_addr_conv_out_mi9;
                                    end
                                 end
                              end
                           end
                           
                        endcase

                     end
                     else begin
                        if (en_0) begin
                           if (en_1) begin
                              if (cycle1_state2) begin
                                 if (drain3) begin
                                 end
                                 else begin
                                    s_reg_1000 <= short_addr_conv_out_mi9;
                                 end
                              end
                              else begin
                                 case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                    7'd001: begin
                                       if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                       end
                                       else begin
                                          s_reg_1000 <= short_addr_conv_out_mi9;
                                       end
                                    end
                                    
                                    default: begin
                                       if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                       end
                                       else begin
                                          s_reg_1000 <= short_addr_conv_out_mi9;
                                       end
                                    end
                                    
                                 endcase

                              end
                           end
                           else begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_1000 <= short_addr_conv_out_mi9;
                              end
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_32bx5i
         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1001
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_1001 <= 32'd0000000000;
                  end
                  
                  5'd01, 5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                        s_reg_1001 <= s_reg_1005[31:0];
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1001 <= bnn_Add_32Ux32U_32U_1_955_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1001 <= bnn_Add_32Ux32U_32U_1_955_out1;
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_1001 <= s_reg_1010;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_1001 <= short_addr_out_fmap_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1001 <= short_addr_out_fmap_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1001 <= short_addr_out_fmap_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_1001 <= short_addr_out_fmap_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_32bx4i
         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1002
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_1002 <= 32'd0000000000;
                  end
                  
                  5'd01: begin
                     s_reg_1002 <= {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1};
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_1002 <= s_reg_1009;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_1002 <= short_addr_in_fmap_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1002 <= short_addr_in_fmap_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1002 <= short_addr_in_fmap_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_1002 <= short_addr_in_fmap_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_32bx4i
         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1003
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_1003 <= 32'd0000000000;
                  end
                  
                  5'd14: begin
                     if (32'd0000000000 != s_reg_1000) begin
                        s_reg_1003 <= {{ 16 {memresp_data[15]}}, memresp_data[15:0]};
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_1003 <= s_reg_1008;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_1003 <= short_addr_kh_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1003 <= short_addr_kh_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1003 <= short_addr_kh_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_1003 <= short_addr_kh_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_1004
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1004 <= bnn_N_Mux_2_2_3_4_62_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1005
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1005 <= bnn_N_Mux_64_2_2_4_63_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1006
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1006 <= bnn_N_Muxb_1_2_18_4_68_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1007
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1007 <= bnn_N_Mux_32_2_1_4_69_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1008
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1008 <= bnn_N_Mux_32_2_1_4_70_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1009
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1009 <= bnn_N_Mux_32_2_1_4_71_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1010
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1010 <= bnn_N_Mux_32_2_1_4_72_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1011
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_1011 <= bnn_N_Mux_32_2_1_4_73_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_3bx5i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_s_reg_1012
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01, 5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                        s_reg_1012 <= 3'd0;
                     end
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1012 <= {1'b0, bnn_N_Mux_2_2_3_1_1420_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1012 <= {1'b0, bnn_N_Mux_2_2_3_1_1420_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1012 <= {2'b00, bnn_GreaterThan_6Sx4S_1U_4_1515_out1};
                        end
                     end
                  end
                  
                  5'd12: begin
                     s_reg_1012 <= bnn_N_Mux_3_2_6_4_4105_out1;
                  end
                  
                  5'd13: begin
                     s_reg_1012 <= bnn_Add_2Ux2U_3U_4_4427_out1;
                  end
                  
               endcase

            end
         end

         // resource: regr_4b
         always @(posedge clk)
          begin :drive_s_reg_1013
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_2) begin
                        case (cycle2_state2) 

                           2'd0, 2'd1: begin
                              if (s_reg_870_stage10) begin
                              end
                              else begin
                                 s_reg_1013 <= bnn_N_Mux_4_2_11_4_83_out1;
                              end
                           end
                           
                        endcase

                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1014
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01, 5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                        s_reg_1014 <= bnn_OrReduction_2U_1U_4_181_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1014 <= bnn_Add_17Sx16S_17S_1_2579_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1014 <= bnn_Add_17Sx16S_17S_1_2579_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1015
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd05, 5'd07: begin
                     s_reg_1015 <= bnn_OrReduction_2U_1U_4_189_out1;
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1015 <= bnn_Add_17Sx16S_17S_1_2606_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1015 <= bnn_Add_17Sx16S_17S_1_2606_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1016
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1016 <= bnn_OrReduction_2U_1U_4_194_out1;
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1016 <= bnn_Add_17Sx16S_17S_1_2633_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1016 <= bnn_Add_17Sx16S_17S_1_2633_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_32bx5i
         // resource: regr_32b
         always @(posedge clk)
          begin :drive_s_reg_1017
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_1017 <= 32'd0000000000;
                  end
                  
                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_1017 <= s_reg_1007;
                        end
                     end
                     else begin
                        s_reg_1017 <= s_reg_1007;
                     end
                  end
                  
                  5'd12: begin
                     s_reg_1017 <= bnn_Add_32Ux10U_32U_1_954_out1;
                  end
                  
                  5'd14: begin
                     if (s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        s_reg_1017 <= 32'd0000000000;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1017 <= {3'b000, bnn_Add_32Ux10U_32U_1_954_out1[28:0]};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1017 <= {3'b000, bnn_Add_32Ux10U_32U_1_954_out1[28:0]};
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_1017 <= s_reg_1007;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_1017 <= short_addr_w_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1017 <= short_addr_w_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_1017 <= short_addr_w_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_1017 <= short_addr_w_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_1018
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_1018_slice <= bnn_N_Mux_4_2_10_4_80_out1_slice;
                        end
                     end
                     else begin
                        s_reg_1018_slice <= bnn_N_Mux_4_2_10_4_80_out1_slice;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_10bx3i
         // resource: regr_10b
         always @(posedge clk)
          begin :drive_s_reg_1019
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                        s_reg_1019 <= 10'd0000;
                     end
                  end
                  
                  5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4] && 32'd0000000000 != s_reg_1005[31:0]) begin
                        s_reg_1019 <= s_reg_1163;
                     end
                  end
                  
                  5'd12: begin
                     s_reg_1019 <= s_reg_1163;
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1019 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4775_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1019 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4775_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_10bx3i
         // resource: regr_10b
         always @(posedge clk)
          begin :drive_s_reg_1020
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        s_reg_1020 <= 10'd0000;
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1020 <= bnn_Add_10Ux1U_10U_4_192_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1020 <= bnn_Add_10Ux1U_10U_4_192_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1020 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4779_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1020 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4779_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_6bx2i
         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1021
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd05, 5'd07: begin
                     s_reg_1021 <= bnn_Mul_30Sx12S_30S_1_191_out1[5:0];
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1021 <= bnn_Add_6Ux6U_6U_1_282_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1021 <= bnn_Add_6Ux6U_6U_1_282_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_3b
         always @(posedge clk)
          begin :drive_s_reg_1022
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd05, 5'd07: begin
                     s_reg_1022 <= bnn_Add_6Sx4S_6S_1_193_out1[2:0];
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1023
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd05, 5'd07: begin
                     s_reg_1023 <= bnn_LessThan_3Ux3U_1U_4_190_out1;
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1023 <= bnn_Add_17Sx16S_17S_1_2660_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1023 <= bnn_Add_17Sx16S_17S_1_2660_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1024
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08, 5'd10: begin
                     s_reg_1024 <= bnn_Not_1U_1U_4_207_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_1024 <= bnn_Not_1U_1U_4_207_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1024 <= bnn_Add_17Sx16S_17S_1_2687_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1024 <= bnn_Add_17Sx16S_17S_1_2687_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx4i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1025
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1025 <= {5'b00000, bnn_Add_7Sx5S_7S_4_195_out1[1:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1025 <= {5'b00000, bnn_Add_7Sx5S_7S_4_195_out1[1:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1025 <= {5'b00000, bnn_N_Mux_2_2_3_1_1394_out1};
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1025 <= {5'b00000, bnn_N_Mux_2_2_3_1_1394_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1025 <= {{ 2 {bnn_Add_7Sx5S_7S_4_195_out1[4]}}, bnn_Add_7Sx5S_7S_4_195_out1[4:0]};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1025 <= bnn_LeftShift_9Ux3U_7U_4_4819_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1025 <= bnn_LeftShift_9Ux3U_7U_4_4819_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_4bx3i
         // resource: regr_4b
         always @(posedge clk)
          begin :drive_s_reg_1026
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1026 <= bnn_Mul_30Sx12S_30S_1_191_out1[3:0];
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1026 <= bnn_Mul_30Sx12S_30S_1_191_out1[3:0];
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1026 <= bnn_Add_4Sx2S_5S_4_1369_out1[3:0];
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1026 <= bnn_Add_4Sx2S_5S_4_1369_out1[3:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1026 <= bnn_Sub_4Ux1U_4S_4_1538_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx3i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1027
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1027 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1027 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1027 <= {bnn_Add_3Sx3S_4S_1_1375_out1[3], bnn_Add_3Sx3S_4S_1_1375_out1};
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1027 <= {bnn_Add_3Sx3S_4S_1_1375_out1[3], bnn_Add_3Sx3S_4S_1_1375_out1};
                        end
                        else begin
                           s_reg_1027 <= bnn_Add_4Sx4S_5S_4_355_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1027 <= bnn_Add_4Sx4S_5S_4_355_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1027 <= bnn_Add_4Sx4S_5S_4_355_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_4bx3i
         // resource: regr_4b
         always @(posedge clk)
          begin :drive_s_reg_1028
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1028 <= bnn_Mul_30Sx12S_30S_1_191_out1[3:0];
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1028 <= bnn_Mul_30Sx12S_30S_1_191_out1[3:0];
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1028 <= bnn_Add_4Sx2S_4S_1_1372_out1;
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1028 <= bnn_Add_4Sx2S_4S_1_1372_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1028 <= bnn_Add_5Sx4S_6S_1_1502_out1[3:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_6bx2i
         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1029
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1029 <= {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_1029 <= {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1029 <= bnn_Add_6Ux6U_6U_1_699_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1029 <= bnn_Add_6Ux6U_6U_1_699_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx3i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1030
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1030 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1030 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1030 <= {3'b000, bnn_N_Mux_2_2_3_4_1455_out1};
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1030 <= {3'b000, bnn_N_Mux_2_2_3_4_1455_out1};
                        end
                        else begin
                           s_reg_1030 <= bnn_Add_4Sx3S_5S_4_463_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1030 <= bnn_Add_4Sx3S_5S_4_463_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1030 <= bnn_Add_4Sx3S_5S_4_463_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_6bx2i
         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1031
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1031 <= {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_1031 <= {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1031 <= bnn_Add_6Ux6U_6U_1_345_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1031 <= bnn_Add_6Ux6U_6U_1_345_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_6bx2i
         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1032
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1032 <= bnn_Add_6Ux6U_6U_1_206_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_1032 <= bnn_Add_6Ux6U_6U_1_206_out1;
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1032 <= bnn_Add_6Ux6U_6U_1_274_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1032 <= bnn_Add_6Ux6U_6U_1_274_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_1033
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08, 5'd10: begin
                     s_reg_1033 <= bnn_Add_2Ux1U_2U_4_208_out1;
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1033 <= bnn_Add_2Ux1U_2U_4_208_out1;
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1033 <= bnn_N_Mux_2_2_3_4_1368_out1;
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1033 <= bnn_N_Mux_2_2_3_4_1368_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1033 <= bnn_Minus_2S_2S_1_1503_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_10bx2i
         // resource: regr_10b
         always @(posedge clk)
          begin :drive_s_reg_1034
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1034 <= s_reg_1020;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1034 <= s_reg_1020;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1034 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4783_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1034 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4783_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx3i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1035
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1035 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1035 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1035 <= bnn_Add_5Sx4S_6S_1_1502_out1[4:0];
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1035 <= bnn_Add_5Sx4S_6S_1_1502_out1[4:0];
                        end
                        else begin
                           s_reg_1035 <= bnn_Add_4Sx4S_5S_4_272_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1035 <= bnn_Add_4Sx4S_5S_4_272_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1035 <= bnn_Add_4Sx4S_5S_4_272_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx3i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1036
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd06, 5'd08: begin
                     s_reg_1036 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_1036 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_1036 <= bnn_Add_6Ux6U_6U_1_409_out1[4:0];
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1036 <= bnn_Add_6Ux6U_6U_1_409_out1[4:0];
                        end
                        else begin
                           s_reg_1036 <= bnn_Add_4Sx2S_5S_4_276_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1036 <= bnn_Add_4Sx2S_5S_4_276_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1036 <= bnn_Add_4Sx2S_5S_4_276_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1037
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1037 <= bnn_GreaterThan_6Sx4S_1U_4_278_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1037 <= bnn_GreaterThan_6Sx4S_1U_4_278_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1037 <= bnn_Add_17Sx16S_17S_1_2824_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1037 <= bnn_Add_17Sx16S_17S_1_2824_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1038
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1038 <= bnn_GreaterThan_6Sx4S_1U_4_286_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1038 <= bnn_GreaterThan_6Sx4S_1U_4_286_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1038 <= bnn_Add_17Sx16S_17S_1_2851_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1038 <= bnn_Add_17Sx16S_17S_1_2851_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1039
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1039 <= bnn_Add_6Ux6U_6U_1_457_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1039 <= bnn_Add_6Ux6U_6U_1_457_out1[4:0];
                        end
                        else begin
                           s_reg_1039 <= bnn_Add_4Sx4S_5S_4_290_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1039 <= bnn_Add_4Sx4S_5S_4_290_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1039 <= bnn_Add_4Sx4S_5S_4_290_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1040
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1040 <= bnn_GreaterThan_6Sx4S_1U_4_294_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1040 <= bnn_GreaterThan_6Sx4S_1U_4_294_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1040 <= bnn_Add_17Sx16S_17S_1_2878_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1040 <= bnn_Add_17Sx16S_17S_1_2878_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1041
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1041 <= {bnn_Add_6Ux6U_6U_1_298_out1[5], bnn_Add_6Ux6U_6U_1_298_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1041 <= {bnn_Add_6Ux6U_6U_1_298_out1[5], bnn_Add_6Ux6U_6U_1_298_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1041 <= bnn_LeftShift_9Ux3U_7U_4_4787_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1041 <= bnn_LeftShift_9Ux3U_7U_4_4787_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1042
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1042 <= bnn_GreaterThan_6Sx4S_1U_4_301_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1042 <= bnn_GreaterThan_6Sx4S_1U_4_301_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1042 <= bnn_Add_17Sx16S_17S_1_2905_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1042 <= bnn_Add_17Sx16S_17S_1_2905_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1043
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1043 <= bnn_Add_6Ux6U_6U_1_699_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1043 <= bnn_Add_6Ux6U_6U_1_699_out1[4:0];
                        end
                        else begin
                           s_reg_1043 <= bnn_Add_4Sx3S_5S_4_304_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1043 <= bnn_Add_4Sx3S_5S_4_304_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1043 <= bnn_Add_4Sx3S_5S_4_304_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1044
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1044 <= bnn_And_1Sx1U_1U_4_305_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1044 <= bnn_And_1Sx1U_1U_4_305_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1044 <= bnn_Add_17Sx16S_17S_1_2714_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1044 <= bnn_Add_17Sx16S_17S_1_2714_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1045
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1045 <= bnn_GreaterThan_6Sx4S_1U_4_308_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1045 <= bnn_GreaterThan_6Sx4S_1U_4_308_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1045 <= bnn_Add_17Sx16S_17S_1_2932_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1045 <= bnn_Add_17Sx16S_17S_1_2932_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1046
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1046 <= {bnn_Add_6Ux6U_6U_1_314_out1[5], bnn_Add_6Ux6U_6U_1_314_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1046 <= {bnn_Add_6Ux6U_6U_1_314_out1[5], bnn_Add_6Ux6U_6U_1_314_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1046 <= bnn_LeftShift_9Ux3U_7U_4_4791_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1046 <= bnn_LeftShift_9Ux3U_7U_4_4791_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1047
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1047 <= bnn_Add_6Ux6U_6U_1_887_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_1047 <= bnn_Add_6Ux6U_6U_1_887_out1[4:0];
                        end
                        else begin
                           s_reg_1047 <= bnn_Add_4Sx4S_5S_4_323_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_1047 <= bnn_Add_4Sx4S_5S_4_323_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_1047 <= bnn_Add_4Sx4S_5S_4_323_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1048
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1048 <= bnn_And_1Sx1U_1U_4_324_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1048 <= bnn_And_1Sx1U_1U_4_324_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1048 <= bnn_Add_17Sx16S_17S_1_2741_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1048 <= bnn_Add_17Sx16S_17S_1_2741_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1049
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1049 <= bnn_GreaterThan_6Sx4S_1U_4_337_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1049 <= bnn_GreaterThan_6Sx4S_1U_4_337_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1049 <= bnn_Add_17Sx16S_17S_1_2957_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1049 <= bnn_Add_17Sx16S_17S_1_2957_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1050
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1050 <= bnn_Or_1Sx1U_1S_4_340_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1050 <= bnn_Or_1Sx1U_1S_4_340_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1050 <= bnn_Add_17Sx16S_17S_1_2769_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1050 <= bnn_Add_17Sx16S_17S_1_2769_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1051
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1051 <= bnn_GreaterThan_6Sx4S_1U_4_347_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1051 <= bnn_GreaterThan_6Sx4S_1U_4_347_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1051 <= bnn_Add_17Sx16S_17S_1_2981_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1051 <= bnn_Add_17Sx16S_17S_1_2981_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1052
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1052 <= bnn_Or_1Sx1U_1S_4_342_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1052 <= bnn_Or_1Sx1U_1S_4_342_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1052 <= bnn_Add_17Sx16S_17S_1_2797_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1052 <= bnn_Add_17Sx16S_17S_1_2797_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1053
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1053 <= bnn_Or_1Sx1U_1S_4_350_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1053 <= bnn_Or_1Sx1U_1S_4_350_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1053 <= bnn_Add_17Sx16S_17S_1_3005_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1053 <= bnn_Add_17Sx16S_17S_1_3005_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1054
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1054 <= bnn_Or_1Sx1U_1S_4_352_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1054 <= bnn_Or_1Sx1U_1S_4_352_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1054 <= bnn_Add_17Sx16S_17S_1_3030_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1054 <= bnn_Add_17Sx16S_17S_1_3030_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1055
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1055 <= bnn_GreaterThan_6Sx4S_1U_4_357_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1055 <= bnn_GreaterThan_6Sx4S_1U_4_357_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1055 <= bnn_Add_17Sx16S_17S_1_3107_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1055 <= bnn_Add_17Sx16S_17S_1_3107_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1056
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1056 <= bnn_Or_1Sx1U_1S_4_360_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1056 <= bnn_Or_1Sx1U_1S_4_360_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1056 <= bnn_Add_17Sx16S_17S_1_3057_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1056 <= bnn_Add_17Sx16S_17S_1_3057_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1057
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1057 <= bnn_Or_1Sx1U_1S_4_362_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1057 <= bnn_Or_1Sx1U_1S_4_362_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1057 <= bnn_Add_17Sx16S_17S_1_3083_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1057 <= bnn_Add_17Sx16S_17S_1_3083_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1058
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1058 <= {bnn_Add_6Ux6U_6U_1_365_out1[5], bnn_Add_6Ux6U_6U_1_365_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1058 <= {bnn_Add_6Ux6U_6U_1_365_out1[5], bnn_Add_6Ux6U_6U_1_365_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1058 <= bnn_LeftShift_9Ux3U_7U_4_4795_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1058 <= bnn_LeftShift_9Ux3U_7U_4_4795_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1059
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1059 <= bnn_LessThanEQ_10Ux33U_1U_4_368_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1059 <= bnn_LessThanEQ_10Ux33U_1U_4_368_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1059 <= bnn_Add_17Sx16S_17S_1_3128_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1059 <= bnn_Add_17Sx16S_17S_1_3128_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1060
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1060 <= bnn_Or_1Sx1U_1S_4_370_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1060 <= bnn_Or_1Sx1U_1S_4_370_out1;
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1060 <= bnn_Add_17Sx16S_17S_1_3146_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1060 <= bnn_Add_17Sx16S_17S_1_3146_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1061
            if (stall0) begin
            end
            else begin
               s_reg_1061 <= bnn_And_1Sx1U_1U_4_374_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1062
            if (stall0) begin
            end
            else begin
               s_reg_1062 <= bnn_GreaterThan_6Sx4S_1U_4_381_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1063
            if (stall0) begin
            end
            else begin
               s_reg_1063 <= bnn_And_1Sx1U_1U_4_386_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1064
            if (stall0) begin
            end
            else begin
               s_reg_1064 <= bnn_OrReduction_10U_1U_4_280_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1065
            if (stall0) begin
            end
            else begin
               s_reg_1065 <= bnn_GreaterThan_6Sx4S_1U_4_503_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1066
            if (stall0) begin
            end
            else begin
               s_reg_1066 <= bnn_And_1Sx1U_1U_4_397_out1;
            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1067
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1067 <= {bnn_Add_6Ux6U_6U_1_407_out1[5], bnn_Add_6Ux6U_6U_1_407_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1067 <= {bnn_Add_6Ux6U_6U_1_407_out1[5], bnn_Add_6Ux6U_6U_1_407_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1067 <= bnn_LeftShift_9Ux3U_7U_4_4799_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1067 <= bnn_LeftShift_9Ux3U_7U_4_4799_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1068
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1068 <= {bnn_Add_6Ux6U_6U_1_409_out1[5], bnn_Add_6Ux6U_6U_1_409_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1068 <= {bnn_Add_6Ux6U_6U_1_409_out1[5], bnn_Add_6Ux6U_6U_1_409_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1068 <= bnn_LeftShift_9Ux3U_7U_4_4803_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1068 <= bnn_LeftShift_9Ux3U_7U_4_4803_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1069
            if (stall0) begin
            end
            else begin
               s_reg_1069 <= bnn_GreaterThan_6Sx4S_1U_4_454_out1;
            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1070
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        s_reg_1070 <= {{ 3 {bnn_LeftShift_2Sx2U_5S_4_75_out1[3]}}, bnn_LeftShift_2Sx2U_5S_4_75_out1[3:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1070 <= bnn_LeftShift_9Ux3U_7U_4_4807_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1070 <= bnn_LeftShift_9Ux3U_7U_4_4807_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1071
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        s_reg_1071 <= bnn_LeftShift_2Sx2U_5S_4_75_out1[3];
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1072
            if (stall0) begin
            end
            else begin
               s_reg_1072 <= bnn_Or_1Sx1U_1S_4_1516_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1073
            if (stall0) begin
            end
            else begin
               s_reg_1073 <= bnn_Or_1Sx1U_1S_4_427_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1074
            if (stall0) begin
            end
            else begin
               s_reg_1074 <= bnn_Or_1Sx1U_1S_4_440_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1075
            if (stall0) begin
            end
            else begin
               s_reg_1075 <= bnn_Or_1Sx1U_1S_4_453_out1;
            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1076
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1076 <= {bnn_Add_6Ux6U_6U_1_457_out1[5], bnn_Add_6Ux6U_6U_1_457_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1076 <= {bnn_Add_6Ux6U_6U_1_457_out1[5], bnn_Add_6Ux6U_6U_1_457_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1076 <= bnn_LeftShift_9Ux3U_7U_4_4811_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1076 <= bnn_LeftShift_9Ux3U_7U_4_4811_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1077
            if (stall0) begin
            end
            else begin
               s_reg_1077 <= s_reg_1076[5];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1078
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        s_reg_1078 <= bnn_OrReduction_2U_1U_4_241_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1079
            if (stall0) begin
            end
            else begin
               s_reg_1079 <= bnn_Or_1Sx1U_1S_4_465_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1080
            if (stall0) begin
            end
            else begin
               s_reg_1080 <= bnn_Or_1Sx1U_1S_4_476_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1081
            if (stall0) begin
            end
            else begin
               s_reg_1081 <= bnn_Or_1Sx1U_1S_4_487_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1082
            if (stall0) begin
            end
            else begin
               s_reg_1082 <= bnn_Or_1Sx1U_1S_4_1517_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1083
            if (stall0) begin
            end
            else begin
               s_reg_1083 <= bnn_Or_1Sx1U_1S_4_498_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1084
            if (stall0) begin
            end
            else begin
               s_reg_1084 <= bnn_Or_1Sx1U_1S_4_1519_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1085
            if (stall0) begin
            end
            else begin
               s_reg_1085 <= bnn_Or_1Sx1U_1S_4_550_out1;
            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1086
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1086 <= bnn_Sub_8Sx2S_8S_4_1520_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1086 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4736_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1086 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4736_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1087
            if (stall0) begin
            end
            else begin
               s_reg_1087 <= s_reg_1029[5];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1088
            if (stall0) begin
            end
            else begin
               s_reg_1088 <= bnn_And_1Sx1U_1U_4_737_out1;
            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1089
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1089 <= bnn_Sub_8Sx2S_8S_4_1522_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1089 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4742_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1089 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4742_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1090
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1090 <= bnn_Sub_8Sx2S_8S_4_1525_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1090 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4751_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1090 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4751_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1091
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1091 <= {{ 2 {bnn_Add_6Ux6U_6U_1_1526_out1[4]}}, bnn_Add_6Ux6U_6U_1_1526_out1[4:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1091 <= {{ 2 {bnn_Add_6Ux6U_6U_1_1526_out1[4]}}, bnn_Add_6Ux6U_6U_1_1526_out1[4:0]};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1091 <= {{ 2 {bnn_Add_6Ux6U_6U_1_1526_out1[4]}}, bnn_Add_6Ux6U_6U_1_1526_out1[4:0]};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1091 <= bnn_LeftShift_9Ux3U_7U_4_4815_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1091 <= bnn_LeftShift_9Ux3U_7U_4_4815_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1092
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1092 <= bnn_Sub_8Sx2S_8S_4_1527_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1092 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4747_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1092 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4747_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1093
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                        if (drain2) begin
                        end
                        else begin
                           s_reg_1093 <= {bnn_Add_6Ux6U_6U_1_887_out1[5], bnn_Add_6Ux6U_6U_1_887_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                        end
                        else begin
                           s_reg_1093 <= {bnn_Add_6Ux6U_6U_1_887_out1[5], bnn_Add_6Ux6U_6U_1_887_out1};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1093 <= bnn_LeftShift_9Ux3U_7U_4_4831_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1093 <= bnn_LeftShift_9Ux3U_7U_4_4831_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1094
            if (stall0) begin
            end
            else begin
               s_reg_1094 <= s_reg_1093[5];
            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1095
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1095 <= {{ 2 {bnn_Add_6Sx4S_6S_1_193_out1[4]}}, bnn_Add_6Sx4S_6S_1_193_out1[4:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1095 <= {{ 2 {bnn_Add_6Sx4S_6S_1_193_out1[4]}}, bnn_Add_6Sx4S_6S_1_193_out1[4:0]};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1095 <= {{ 2 {bnn_Add_6Sx4S_6S_1_193_out1[4]}}, bnn_Add_6Sx4S_6S_1_193_out1[4:0]};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1095 <= bnn_LeftShift_9Ux3U_7U_4_4823_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1095 <= bnn_LeftShift_9Ux3U_7U_4_4823_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1096
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1096 <= bnn_Sub_8Sx2S_8S_4_1529_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1096 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4767_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1096 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4767_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1097
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1097 <= {{ 2 {bnn_Add_5Sx4S_6S_1_212_out1[4]}}, bnn_Add_5Sx4S_6S_1_212_out1[4:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1097 <= {{ 2 {bnn_Add_5Sx4S_6S_1_212_out1[4]}}, bnn_Add_5Sx4S_6S_1_212_out1[4:0]};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1097 <= {{ 2 {bnn_Add_5Sx4S_6S_1_212_out1[4]}}, bnn_Add_5Sx4S_6S_1_212_out1[4:0]};
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1097 <= bnn_LeftShift_9Ux3U_7U_4_4827_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1097 <= bnn_LeftShift_9Ux3U_7U_4_4827_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1098
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1098 <= bnn_Sub_8Sx2S_8S_4_1531_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1098 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4771_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1098 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4771_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1099
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1099 <= {3'b000, bnn_N_Mux_2_2_3_1_1407_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1099 <= {3'b000, bnn_N_Mux_2_2_3_1_1407_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1099 <= bnn_Add_5Sx4S_6S_1_213_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1100
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1100 <= bnn_Sub_8Sx2S_8S_4_1533_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1100 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4755_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1100 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4755_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1101
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1101 <= {{ 2 {bnn_Add_5Sx4S_6S_1_214_out1[4]}}, bnn_Add_5Sx4S_6S_1_214_out1[4:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1101 <= bnn_LeftShift_9Ux3U_7U_4_4839_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1101 <= bnn_LeftShift_9Ux3U_7U_4_4839_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1102
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1102 <= {{ 2 {bnn_Add_5Sx4S_6S_1_215_out1[4]}}, bnn_Add_5Sx4S_6S_1_215_out1[4:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1102 <= bnn_LeftShift_9Ux3U_7U_4_4843_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1102 <= bnn_LeftShift_9Ux3U_7U_4_4843_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1103
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1103 <= bnn_Sub_8Sx2S_8S_4_1536_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1103 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4759_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1103 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4759_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1104
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1104 <= {{ 2 {bnn_Add_5Sx4S_6S_1_216_out1[4]}}, bnn_Add_5Sx4S_6S_1_216_out1[4:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1104 <= bnn_LeftShift_9Ux3U_7U_4_4850_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1104 <= bnn_LeftShift_9Ux3U_7U_4_4850_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_8bx2i
         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1105
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1105 <= bnn_Sub_8Sx2S_8S_4_1540_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1105 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4763_out1};
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1105 <= {1'b0, bnn_LeftShift_9Ux3U_7U_4_4763_out1};
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1106
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1106 <= {{ 2 {bnn_Add_5Sx4S_6S_1_1542_out1[4]}}, bnn_Add_5Sx4S_6S_1_1542_out1[4:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1106 <= bnn_LeftShift_9Ux3U_7U_4_4852_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1106 <= bnn_LeftShift_9Ux3U_7U_4_4852_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx2i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_1107
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd11: begin
                     if (cycle1_state) begin
                     end
                     else begin
                        s_reg_1107 <= {{ 2 {bnn_Add_7Sx4S_7S_1_227_out1[4]}}, bnn_Add_7Sx4S_7S_1_227_out1[4:0]};
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_1107 <= bnn_LeftShift_9Ux3U_7U_4_4854_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_1107 <= bnn_LeftShift_9Ux3U_7U_4_4854_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1108
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1108 <= {3'b000, bnn_N_Mux_2_2_3_4_3724_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1108 <= {3'b000, bnn_N_Mux_2_2_3_4_3724_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1108 <= bnn_Add_5Sx4S_6S_4_1552_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1109
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1109 <= {3'b000, bnn_N_Mux_2_2_3_4_3774_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1109 <= {3'b000, bnn_N_Mux_2_2_3_4_3774_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1109 <= bnn_Add_5Sx4S_6S_4_1556_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1110
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1110 <= {3'b000, bnn_N_Mux_2_2_3_4_1472_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1110 <= {3'b000, bnn_N_Mux_2_2_3_4_1472_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1110 <= bnn_Add_5Sx4S_6S_4_1565_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1111
            if (stall0) begin
            end
            else begin
               s_reg_1111 <= bnn_And_1Sx1U_1U_4_952_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1112
            if (stall0) begin
            end
            else begin
               s_reg_1112 <= bnn_LessThan_10Ux32U_1U_4_1576_out1;
            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1113
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1113 <= {3'b000, bnn_N_Mux_2_2_3_1_1293_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1113 <= {3'b000, bnn_N_Mux_2_2_3_1_1293_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1113 <= bnn_Add_4Sx2S_5S_1_1034_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1114
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1114 <= {3'b000, bnn_N_Mux_2_2_3_4_3849_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1114 <= {3'b000, bnn_N_Mux_2_2_3_4_3849_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1114 <= bnn_Add_4Sx2S_5S_1_1037_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1115
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1115 <= {3'b000, bnn_N_Mux_2_2_3_1_1384_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1115 <= {3'b000, bnn_N_Mux_2_2_3_1_1384_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1115 <= bnn_Add_4Sx2S_5S_1_1057_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1116
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1116 <= {3'b000, bnn_N_Mux_2_2_3_1_1294_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1116 <= {3'b000, bnn_N_Mux_2_2_3_1_1294_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1116 <= bnn_Add_4Sx2S_5S_1_1075_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1117
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1117 <= {3'b000, bnn_N_Mux_2_2_3_4_4054_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1117 <= {3'b000, bnn_N_Mux_2_2_3_4_4054_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1117 <= bnn_Add_4Sx2S_5S_1_1092_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1118
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1118 <= {3'b000, bnn_N_Mux_2_2_3_4_1285_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1118 <= {3'b000, bnn_N_Mux_2_2_3_4_1285_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1118 <= bnn_Add_4Sx2S_5S_4_1109_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1119
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1119 <= {3'b000, bnn_N_Mux_2_2_3_4_1286_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1119 <= {3'b000, bnn_N_Mux_2_2_3_4_1286_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1119 <= bnn_Add_4Sx2S_5S_1_1125_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1120
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1120 <= {3'b000, bnn_N_Mux_2_2_3_1_4076_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1120 <= {3'b000, bnn_N_Mux_2_2_3_1_4076_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1120 <= bnn_Add_4Sx2S_5S_1_1137_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1121
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1121 <= {3'b000, bnn_N_Mux_2_2_3_1_4078_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1121 <= {3'b000, bnn_N_Mux_2_2_3_1_4078_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1121 <= bnn_Add_4Sx2S_5S_1_1154_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1122
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1122 <= {3'b000, bnn_N_Mux_2_2_3_1_4080_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1122 <= {3'b000, bnn_N_Mux_2_2_3_1_4080_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1122 <= bnn_Add_4Sx2S_5S_1_1173_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1123
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1123 <= {3'b000, bnn_N_Mux_2_2_3_1_1371_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1123 <= {3'b000, bnn_N_Mux_2_2_3_1_1371_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1123 <= bnn_Add_4Sx2S_5S_1_1193_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx2i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1124
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1124 <= {3'b000, bnn_N_Mux_2_2_3_1_1374_out1};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1124 <= {3'b000, bnn_N_Mux_2_2_3_1_1374_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1124 <= bnn_Add_4Sx2S_5S_1_1211_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1125
            if (stall0) begin
            end
            else begin
               s_reg_1125 <= bnn_Add_4Sx2S_5S_1_1228_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1126
            if (stall0) begin
            end
            else begin
               s_reg_1126 <= bnn_Add_4Sx2S_5S_1_1245_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1127
            if (stall0) begin
            end
            else begin
               s_reg_1127 <= bnn_Add_4Sx2S_5S_1_1261_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1128
            if (stall0) begin
            end
            else begin
               s_reg_1128 <= bnn_Add_4Sx2S_5S_1_1269_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1129
            if (stall0) begin
            end
            else begin
               s_reg_1129 <= bnn_Add_4Sx2S_5S_1_1280_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1130
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1130 <= bnn_Add_5Sx4S_6S_4_1313_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1130 <= bnn_Add_5Sx4S_6S_4_1313_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1130 <= bnn_Add_5Sx4S_6S_4_1313_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1131
            if (stall0) begin
            end
            else begin
               s_reg_1131 <= bnn_Add_4Sx2S_5S_1_1340_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1132
            if (stall0) begin
            end
            else begin
               s_reg_1132 <= bnn_Add_4Sx2S_5S_4_1355_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1133
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1133 <= bnn_Add_4Sx2S_5S_4_1367_out1;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1133 <= bnn_Add_4Sx2S_5S_4_1367_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1133 <= bnn_Add_4Sx2S_5S_4_1367_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1134
            if (stall0) begin
            end
            else begin
               s_reg_1134 <= bnn_Add_4Sx2S_5S_4_1378_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1135
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1135 <= bnn_Add_5Sx4S_6S_1_1389_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1135 <= bnn_Add_5Sx4S_6S_1_1389_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1135 <= bnn_Add_5Sx4S_6S_1_1389_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1136
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1136 <= bnn_Add_5Sx4S_6S_1_1400_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1136 <= bnn_Add_5Sx4S_6S_1_1400_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1136 <= bnn_Add_5Sx4S_6S_1_1400_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1137
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1137 <= bnn_Add_5Sx4S_6S_4_1426_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1137 <= bnn_Add_5Sx4S_6S_4_1426_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1137 <= bnn_Add_5Sx4S_6S_4_1426_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_16bx2i
         // resource: regr_16b
         always @(posedge clk)
          begin :drive_s_reg_1138
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1138 <= {{ 11 {bnn_Add_5Sx4S_6S_1_1443_out1[4]}}, bnn_Add_5Sx4S_6S_1_1443_out1[4:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1138 <= {{ 11 {bnn_Add_5Sx4S_6S_1_1443_out1[4]}}, bnn_Add_5Sx4S_6S_1_1443_out1[4:0]};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1138 <= {{ 11 {bnn_Add_5Sx4S_6S_1_1443_out1[4]}}, bnn_Add_5Sx4S_6S_1_1443_out1[4:0]};
                        end
                     end
                  end
                  
                  5'd14: begin
                     if (32'd0000000000 != s_reg_1000) begin
                        s_reg_1138 <= memresp_data[31:16];
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1139
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1139 <= bnn_Add_5Sx4S_6S_1_1460_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1139 <= bnn_Add_5Sx4S_6S_1_1460_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1139 <= bnn_Add_5Sx4S_6S_1_1460_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1140
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1140 <= bnn_Add_5Sx4S_6S_1_1475_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1140 <= bnn_Add_5Sx4S_6S_1_1475_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1140 <= bnn_Add_5Sx4S_6S_1_1475_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1141
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1141 <= bnn_Add_5Sx4S_6S_1_1487_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1141 <= bnn_Add_5Sx4S_6S_1_1487_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1141 <= bnn_Add_5Sx4S_6S_1_1487_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1142
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1142 <= bnn_Add_5Sx4S_6S_1_1496_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1142 <= bnn_Add_5Sx4S_6S_1_1496_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1142 <= bnn_Add_5Sx4S_6S_1_1496_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1143
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_1143 <= bnn_Add_5Sx4S_6S_1_1501_out1[4:0];
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_1143 <= bnn_Add_5Sx4S_6S_1_1501_out1[4:0];
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_1143 <= bnn_Add_5Sx4S_6S_1_1501_out1[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1144
            if (stall0) begin
            end
            else begin
               s_reg_1144 <= bnn_N_Mux_64_2_2_1_4563_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1145
            if (stall0) begin
            end
            else begin
               s_reg_1145 <= bnn_N_Mux_64_2_2_1_4572_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1146
            if (stall0) begin
            end
            else begin
               s_reg_1146 <= bnn_N_Mux_64_2_2_1_4581_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1147
            if (stall0) begin
            end
            else begin
               s_reg_1147 <= bnn_N_Mux_64_2_2_1_4590_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1148
            if (stall0) begin
            end
            else begin
               s_reg_1148 <= bnn_N_Mux_64_2_2_1_4599_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1149
            if (stall0) begin
            end
            else begin
               s_reg_1149 <= bnn_N_Mux_64_2_2_1_4608_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1150
            if (stall0) begin
            end
            else begin
               s_reg_1150 <= bnn_N_Mux_64_2_2_1_4617_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1151
            if (stall0) begin
            end
            else begin
               s_reg_1151 <= bnn_N_Mux_64_2_2_1_4626_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1152
            if (stall0) begin
            end
            else begin
               s_reg_1152 <= bnn_N_Mux_64_2_2_1_4635_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1153
            if (stall0) begin
            end
            else begin
               s_reg_1153 <= bnn_N_Mux_64_2_2_1_4644_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1154
            if (stall0) begin
            end
            else begin
               s_reg_1154 <= bnn_N_Mux_64_2_2_1_4653_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1155
            if (stall0) begin
            end
            else begin
               s_reg_1155 <= bnn_N_Mux_64_2_2_1_4662_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1156
            if (stall0) begin
            end
            else begin
               s_reg_1156 <= bnn_N_Mux_64_2_2_1_4671_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1157
            if (stall0) begin
            end
            else begin
               s_reg_1157 <= bnn_N_Mux_64_2_2_1_4680_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1158
            if (stall0) begin
            end
            else begin
               s_reg_1158 <= bnn_N_Mux_64_2_2_1_4689_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1159
            if (stall0) begin
            end
            else begin
               s_reg_1159 <= bnn_N_Mux_64_2_2_1_4698_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1160
            if (stall0) begin
            end
            else begin
               s_reg_1160 <= bnn_N_Mux_64_2_2_1_4707_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1161
            if (stall0) begin
            end
            else begin
               s_reg_1161 <= bnn_N_Mux_64_2_2_1_4716_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1162
            if (stall0) begin
            end
            else begin
               s_reg_1162 <= bnn_N_Mux_64_2_2_1_4725_out1;
            end
         end

         // resource: mux_10bx4i
         // resource: regr_10b
         always @(posedge clk)
          begin :drive_s_reg_1163
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     s_reg_1163 <= 10'd0000;
                  end
                  
                  5'd05, 5'd07: begin
                     s_reg_1163 <= bnn_Add_10Ux1U_10U_4_192_out1;
                  end
                  
                  5'd14: begin
                     if (32'd0000000000 == s_reg_1000) begin
                        s_reg_1163 <= 10'd0000;
                     end
                  end
                  
                  5'd15: begin
                     if (!cycle3_state && !s_reg_1044_stage2) begin
                        if (drain1) begin
                           s_reg_1163 <= 10'd0000;
                        end
                        else begin
                           s_reg_1163 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4729_out1};
                        end
                     end
                     else begin
                        if (cycle1_state0) begin
                           if (drain1) begin
                           end
                           else begin
                              s_reg_1163 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4729_out1};
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                           end
                           else begin
                              s_reg_1163 <= {3'b000, bnn_LeftShift_9Ux3U_7U_4_4729_out1};
                           end
                        end
                     end
                  end
                  
                  5'd16: begin
                     if (!cycle2_state1 && !s_reg_907) begin
                        s_reg_1163 <= 10'd0000;
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                        if (s_reg_907) begin
                        end
                        else begin
                           s_reg_1163 <= 10'd0000;
                        end
                     end
                     else begin
                        s_reg_1163 <= {3'b000, bnn_Add_7Sx5S_7S_4_195_out1};
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1164
            if (stall0) begin
            end
            else begin
               s_reg_1164 <= bnn_N_Mux_64_2_2_1_4733_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1165
            if (stall0) begin
            end
            else begin
               s_reg_1165 <= bnn_N_Mux_64_2_2_1_4740_out1;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_1166
            if (stall0) begin
            end
            else begin
               s_reg_1166 <= bnn_N_Mux_64_2_2_1_4746_out1;
            end
         end

         // resource: mux_1bx5i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_870
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_870 <= 1'b1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_870 <= bnn_OrReduction_2U_1U_4_3548_out1;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_870 <= bnn_OrReduction_2U_1U_4_3548_out1;
                        end
                        else begin
                           s_reg_870 <= bnn_And_1Sx1U_1U_4_315_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_870 <= bnn_And_1Sx1U_1U_4_315_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_870 <= bnn_And_1Sx1U_1U_4_315_out1;
                           end
                        end
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_870 <= bnn_Add_17Sx16S_17S_1_3546_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_870 <= bnn_Add_17Sx16S_17S_1_3546_out1[16];
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_870 <= 1'b1;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_870 <= short_popped_go_0_u0_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_870 <= short_popped_go_0_u0_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_870 <= short_popped_go_0_u0_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_870 <= short_popped_go_0_u0_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_5bx6i
         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_871
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01, 5'd02: begin
                     s_reg_871 <= bnn_Add_5Sx4S_6S_1_180_out1[4:0];
                  end
                  
                  5'd06, 5'd08: begin
                     s_reg_871 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  
                  5'd09: begin
                     if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     end
                     else begin
                        if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                           s_reg_871 <= {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                        end
                        else begin
                           if (32'd0000000000 == s_reg_1000) begin
                              s_reg_871 <= bnn_Add_5Sx4S_6S_1_180_out1[4:0];
                           end
                        end
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        if (drain2) begin
                           s_reg_871 <= bnn_Add_5Sx4S_6S_1_180_out1[4:0];
                        end
                        else begin
                           s_reg_871 <= bnn_LeftShift_2Sx2U_5S_4_75_out1;
                        end
                     end
                     else begin
                        if (cycle1_state) begin
                           if (drain2) begin
                           end
                           else begin
                              s_reg_871 <= bnn_LeftShift_2Sx2U_5S_4_75_out1;
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_2_out1) begin
                           end
                           else begin
                              s_reg_871 <= bnn_LeftShift_2Sx2U_5S_4_75_out1;
                           end
                        end
                     end
                  end
                  
                  5'd14: begin
                     s_reg_871 <= 5'd00;
                  end
                  
                  5'd15: begin
                     if (!cycle3_state && !s_reg_1044_stage2) begin
                        if (drain1) begin
                           s_reg_871 <= 5'd00;
                        end
                        else begin
                           s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                        end
                     end
                     else begin
                        if (cycle1_state0) begin
                           if (drain1) begin
                           end
                           else begin
                              s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                           end
                           else begin
                              s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                           end
                        end
                     end
                  end
                  
                  5'd16: begin
                     if (!cycle2_state1 && !s_reg_907) begin
                        if (drain) begin
                           s_reg_871 <= 5'd00;
                        end
                        else begin
                           s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                        end
                     end
                     else begin
                        if (cycle1_state1) begin
                           if (drain) begin
                           end
                           else begin
                              s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                           end
                        end
                        else begin
                           if (bnn_Equal_1Ux1U_1U_1_1_4_out1) begin
                           end
                           else begin
                              s_reg_871 <= bnn_Add_6Sx4S_6S_1_193_out1[4:0];
                           end
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                        if (s_reg_907) begin
                        end
                        else begin
                           s_reg_871 <= s_reg_886[4:0];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_872
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_872 <= 2'd0;
                  end
                  
                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_872 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_872 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_872 <= bnn_N_Mux_2_2_3_1_3071_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_872 <= bnn_N_Mux_2_2_3_1_3071_out1;
                           end
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_872 <= s_reg_1004;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_872 <= short_width_mode_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_872 <= short_width_mode_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_872 <= short_width_mode_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_872 <= short_width_mode_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_873
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_873 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_873 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_873 <= bnn_N_Mux_2_2_3_1_3093_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_873 <= bnn_N_Mux_2_2_3_1_3093_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx6i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_874
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_874 <= 7'd000;
                        end
                     end
                     else begin
                        s_reg_874 <= 7'd000;
                     end
                  end
                  
                  5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_874 <= {{ 5 {s_reg_874[1]}}, s_reg_874[1:0]};
                        end
                     end
                     else begin
                        s_reg_874 <= {{ 5 {s_reg_874[1]}}, s_reg_874[1:0]};
                     end
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_874 <= {{ 5 {s_reg_874[1]}}, s_reg_874[1:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_874 <= {{ 5 {bnn_N_Mux_2_2_3_1_1831_out1[1]}}, bnn_N_Mux_2_2_3_1_1831_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (s_reg_1000 != 32'd0000000000 && !s_reg_1071) begin
                              s_reg_874 <= {{ 2 {bnn_Add_5Sx3S_5S_1_209_out1[4]}}, bnn_Add_5Sx3S_5S_1_209_out1};
                           end
                           else begin
                              s_reg_874 <= {{ 5 {Bline_buffer_1_mi61[1]}}, Bline_buffer_1_mi61};
                           end
                        end
                     end
                  end
                  
                  5'd12: begin
                     s_reg_874 <= {{ 5 {s_reg_874[1]}}, s_reg_874[1:0]};
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_874 <= bnn_LeftShift_9Ux3U_7U_4_4847_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_874 <= bnn_LeftShift_9Ux3U_7U_4_4847_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_875
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_875 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_875 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_875 <= bnn_N_Mux_2_2_3_1_1846_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_875 <= Bline_buffer_2_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_876
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_876 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_876 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_876 <= {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_876 <= Bline_buffer_11_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_877
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_877 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_877 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_877 <= {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_877 <= Bline_buffer_12_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_878
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_878 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_878 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_878 <= bnn_N_Mux_2_2_3_1_3114_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_878 <= bnn_N_Mux_2_2_3_1_3114_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_879
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_879 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_879 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_879 <= bnn_N_Mux_2_2_3_1_1933_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (s_reg_1004 == 2'd1 && s_reg_1000 != 32'd0000000000) begin
                              s_reg_879 <= bnn_N_Mux_3_2_6_4_957_out1_slice;
                           end
                           else begin
                              s_reg_879 <= Bline_buffer_31_mi61;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_880
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_880 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_880 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_880 <= bnn_N_Mux_2_2_3_1_1944_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_880 <= Bline_buffer_32_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_881
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_881 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_881 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_881 <= bnn_N_Mux_2_2_3_1_1857_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_881 <= Bline_buffer_3_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_882
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_882 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_882 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_882 <= {bnn_N_Mux_64_2_2_1_1636_out1[34], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_882 <= Bline_buffer_13_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_883
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_883 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_883 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_883 <= bnn_N_Mux_3_2_6_4_2178_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_883 <= bnn_N_Mux_3_2_6_4_959_out1_slice;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_884
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_884 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_884 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_884 <= bnn_N_Mux_2_2_3_1_3133_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_884 <= bnn_N_Mux_2_2_3_1_3133_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_885
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_885 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_885 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_885 <= bnn_N_Mux_2_2_3_1_1955_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_885 <= Bline_buffer_33_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_7bx6i
         // resource: regr_7b
         always @(posedge clk)
          begin :drive_s_reg_886
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_886 <= 7'd000;
                        end
                     end
                     else begin
                        s_reg_886 <= 7'd000;
                     end
                  end
                  
                  5'd02: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_886 <= {{ 5 {s_reg_886[1]}}, s_reg_886[1:0]};
                        end
                     end
                     else begin
                        s_reg_886 <= {{ 5 {s_reg_886[1]}}, s_reg_886[1:0]};
                     end
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 == s_reg_1000)) begin
                        s_reg_886 <= {{ 5 {s_reg_886[1]}}, s_reg_886[1:0]};
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_886 <= {{ 5 {bnn_N_Mux_2_2_3_1_3216_out1[1]}}, bnn_N_Mux_2_2_3_1_3216_out1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (s_reg_1000 != 32'd0000000000 && !s_reg_1076[5]) begin
                              s_reg_886 <= {{ 2 {bnn_Add_5Sx4S_6S_1_180_out1[4]}}, bnn_Add_5Sx4S_6S_1_180_out1[4:0]};
                           end
                           else begin
                              if (cycle2_state) begin
                                 s_reg_886 <= {{ 5 {s_reg_886[1]}}, s_reg_886[1:0]};
                              end
                              else begin
                                 s_reg_886 <= {{ 5 {bnn_N_Mux_2_2_3_1_3216_out1[1]}}, bnn_N_Mux_2_2_3_1_3216_out1};
                              end
                           end
                        end
                     end
                  end
                  
                  5'd12: begin
                     s_reg_886 <= {{ 5 {s_reg_886[1]}}, s_reg_886[1:0]};
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_886 <= bnn_LeftShift_9Ux3U_7U_4_4835_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_886 <= bnn_LeftShift_9Ux3U_7U_4_4835_out1;
                        end
                     end
                  end
                  
                  5'd17: begin
                     s_reg_886 <= {2'b00, bnn_Add_5Sx4S_6S_1_180_out1[4:0]};
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_887
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_887 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_887 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_887 <= bnn_N_Mux_3_2_6_4_1922_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_887 <= bnn_Minus_2S_2S_4_960_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_888
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_888 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_888 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_888 <= bnn_N_Mux_2_2_3_1_1868_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_888 <= Bline_buffer_4_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_889
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_889 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_889 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_889 <= {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_889 <= Bline_buffer_14_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_890
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_890 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_890 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_890 <= bnn_N_Mux_2_2_3_1_3151_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_890 <= bnn_N_Mux_2_2_3_1_3151_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_891
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_891 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_891 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_891 <= bnn_N_Mux_2_2_3_1_2176_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_891 <= Bline_buffer_30_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_892
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_892 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_892 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_892 <= bnn_N_Mux_2_2_3_1_1966_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_892 <= Bline_buffer_34_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_893
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_893 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_893 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_893 <= {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_893 <= Bline_buffer_41_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_894
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_894 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_894 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_894 <= bnn_N_Mux_2_2_3_1_3203_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_894 <= bnn_N_Mux_2_2_3_1_3203_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_895
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_895 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_895 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_895 <= bnn_N_Mux_2_2_3_1_3229_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_895 <= bnn_N_Mux_2_2_3_1_3229_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_896
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_896 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_896 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_896 <= bnn_N_Mux_2_2_3_1_2021_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_896 <= Bline_buffer_61_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_64bx5i
         // resource: regr_64b
         always @(posedge clk)
          begin :drive_s_reg_897
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00, 5'd01: begin
                     s_reg_897 <= 64'd00000000000000000000;
                  end
                  
                  5'd08: begin
                     s_reg_897 <= memresp_data[63:0];
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_897 <= bnn_And_64Sx64S_64S_1_4562_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_897 <= bnn_And_64Sx64S_64S_1_4562_out1;
                        end
                     end
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_897 <= s_reg_1005;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_897 <= short_n_inputs_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_897 <= short_n_inputs_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_897 <= short_n_inputs_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_897 <= short_n_inputs_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_898
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_898 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_898 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_898 <= bnn_N_Mux_2_2_3_1_1879_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_898 <= Bline_buffer_5_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_899
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_899 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_899 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_899 <= {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_899 <= Bline_buffer_15_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_900
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_900 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_900 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_900 <= bnn_N_Mux_2_2_3_1_3168_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_900 <= bnn_N_Mux_2_2_3_1_3168_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_901
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_901 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_901 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_901 <= bnn_N_Mux_2_2_3_1_1977_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_901 <= Bline_buffer_35_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_902
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_902 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_902 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_902 <= bnn_N_Mux_3_2_6_4_1638_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_902 <= Bline_buffer_40_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_903
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_903 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_903 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_903 <= {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_903 <= Bline_buffer_42_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_904
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_904 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_904 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_904 <= bnn_N_Mux_2_2_3_1_3243_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_904 <= bnn_N_Mux_2_2_3_1_3243_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_905
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_905 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_905 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_905 <= bnn_N_Mux_2_2_3_1_2208_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_905 <= Bline_buffer_60_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_906
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_906 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_906 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_906 <= bnn_N_Mux_2_2_3_1_2038_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_906 <= Bline_buffer_62_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx7i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_907
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     s_reg_907 <= 1'b0;
                  end
                  
                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_907 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_907 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_907 <= bnn_N_Muxb_1_2_18_4_230_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_907 <= bnn_N_Muxb_1_2_18_4_230_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_907 <= bnn_Equal_2Ux2U_1U_4_4460_out1;
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_907 <= bnn_Equal_2Ux2U_1U_4_4460_out1;
                        end
                     end
                  end
                  
                  5'd16: begin
                     if (cycle1_state1) begin
                     end
                     else begin
                        s_reg_907 <= bnn_LessThan_5Ux32U_1U_4_5204_out1;
                     end
                  end
                  
                  5'd17: begin
                     s_reg_907 <= bnn_Add_5Sx4S_6S_1_180_out1[4];
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        s_reg_907 <= s_reg_1006;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              if (drain3) begin
                              end
                              else begin
                                 s_reg_907 <= short_do_max_pool_mi9;
                              end
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_907 <= short_do_max_pool_mi9;
                                    end
                                 end
                                 
                                 default: begin
                                    if (bnn_Equal_1Ux1U_1U_1_1_out1) begin
                                    end
                                    else begin
                                       s_reg_907 <= short_do_max_pool_mi9;
                                    end
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           if (drain3) begin
                           end
                           else begin
                              s_reg_907 <= short_do_max_pool_mi9;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_908
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_908 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_908 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_908 <= bnn_N_Muxb_1_2_18_4_229_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_908 <= bnn_N_Muxb_1_2_18_4_229_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_908 <= bnn_Add_17Sx16S_17S_1_3547_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_908 <= bnn_Add_17Sx16S_17S_1_3547_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_909
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_909 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_909 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_909 <= bnn_N_Mux_2_2_3_1_1890_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_909 <= Bline_buffer_6_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_910
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_910 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_910 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_910 <= {bnn_N_Mux_64_2_2_1_1636_out1[37], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_910 <= Bline_buffer_16_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_911
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_911 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_911 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_911 <= bnn_N_Mux_2_2_3_1_3184_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_911 <= bnn_N_Mux_2_2_3_1_3184_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_912
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_912 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_912 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_912 <= bnn_N_Mux_2_2_3_1_1988_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_912 <= Bline_buffer_36_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_913
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_913 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_913 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_913 <= {bnn_N_Mux_64_2_2_1_1636_out1[42], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_913 <= Bline_buffer_43_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_914
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_914 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_914 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_914 <= bnn_N_Mux_2_2_3_1_3258_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_914 <= bnn_N_Mux_2_2_3_1_3258_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_915
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_915 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_915 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_915 <= bnn_N_Mux_2_2_3_1_2055_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_915 <= Bline_buffer_63_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_916
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_916 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_916 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_916 <= bnn_N_Muxb_1_2_18_4_231_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_916 <= bnn_N_Muxb_1_2_18_4_231_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_916 <= bnn_Add_17Sx16S_17S_1_2390_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_916 <= bnn_Add_17Sx16S_17S_1_2390_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_917
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_917 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_917 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_917 <= bnn_N_Mux_2_2_3_1_1901_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_917 <= Bline_buffer_7_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_918
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_918 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_918 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_918 <= {bnn_N_Mux_64_2_2_1_1636_out1[38], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_918 <= Bline_buffer_17_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_919
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_919 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_919 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_919 <= bnn_N_Mux_2_2_3_4_3200_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_919 <= bnn_N_Mux_2_2_3_4_3200_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_920
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_920 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_920 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_920 <= bnn_N_Mux_2_2_3_1_1999_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_920 <= Bline_buffer_37_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_921
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_921 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_921 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_921 <= {bnn_N_Mux_64_2_2_1_1636_out1[43], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_921 <= Bline_buffer_44_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_922
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_922 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_922 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_922 <= bnn_N_Mux_2_2_3_1_3274_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_922 <= bnn_N_Mux_2_2_3_1_3274_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_923
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_923 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_923 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_923 <= bnn_N_Mux_2_2_3_1_2072_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_923 <= Bline_buffer_64_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_924
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_924 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_924 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_924 <= bnn_N_Muxb_1_2_18_4_232_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_924 <= bnn_N_Muxb_1_2_18_4_232_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_924 <= bnn_Add_17Sx16S_17S_1_2417_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_924 <= bnn_Add_17Sx16S_17S_1_2417_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_925
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_925 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_925 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_925 <= bnn_N_Mux_2_2_3_1_1912_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_925 <= Bline_buffer_8_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_926
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_926 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_926 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_926 <= {bnn_N_Mux_64_2_2_1_1636_out1[39], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_926 <= Bline_buffer_18_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_927
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_927 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_927 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_927 <= bnn_N_Mux_2_2_3_1_3215_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_927 <= bnn_N_Mux_2_2_3_1_3215_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_928
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_928 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_928 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_928 <= bnn_N_Mux_2_2_3_1_2010_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_928 <= Bline_buffer_38_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_929
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_929 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_929 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_929 <= {bnn_N_Mux_64_2_2_1_1636_out1[44], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_929 <= Bline_buffer_45_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_930
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_930 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_930 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_930 <= bnn_N_Mux_2_2_3_1_3290_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_930 <= bnn_N_Mux_2_2_3_1_3290_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_931
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_931 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_931 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_931 <= bnn_N_Mux_2_2_3_1_2089_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_931 <= Bline_buffer_65_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_932
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_932 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_932 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_932 <= bnn_N_Muxb_1_2_18_4_233_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_932 <= bnn_N_Muxb_1_2_18_4_233_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_932 <= bnn_Add_17Sx16S_17S_1_2444_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_932 <= bnn_Add_17Sx16S_17S_1_2444_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_933
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_933 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_933 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_933 <= bnn_N_Mux_2_2_3_1_2164_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_933 <= Bline_buffer_9_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_934
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_934 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_934 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_934 <= bnn_N_Mux_3_2_6_4_1637_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_934 <= Bline_buffer_19_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_935
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_935 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_935 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_935 <= bnn_N_Mux_2_2_3_1_2190_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_935 <= Bline_buffer_39_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_936
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_936 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_936 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_936 <= {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_936 <= Bline_buffer_46_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_937
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_937 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_937 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_937 <= bnn_N_Mux_2_2_3_1_3306_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_937 <= bnn_N_Mux_2_2_3_1_3306_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_938
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_938 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_938 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_938 <= bnn_N_Mux_2_2_3_1_2106_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_938 <= Bline_buffer_66_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_939
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_939 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_939 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_939 <= bnn_N_Muxb_1_2_18_4_234_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_939 <= bnn_N_Muxb_1_2_18_4_234_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_939 <= bnn_Add_17Sx16S_17S_1_2471_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_939 <= bnn_Add_17Sx16S_17S_1_2471_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_940
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_940 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_940 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_940 <= {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_940 <= Bline_buffer_47_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_941
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_941 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_941 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_941 <= bnn_N_Mux_2_2_3_1_3322_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_941 <= bnn_N_Mux_2_2_3_1_3322_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_942
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_942 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_942 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_942 <= bnn_N_Mux_2_2_3_1_2123_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_942 <= Bline_buffer_67_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_943
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_943 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_943 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_943 <= bnn_N_Mux_2_2_3_4_3325_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_943 <= bnn_N_Mux_2_2_3_4_3325_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_944
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_944 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_944 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_944 <= bnn_N_Muxb_1_2_18_4_235_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_944 <= bnn_N_Muxb_1_2_18_4_235_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_944 <= bnn_Add_17Sx16S_17S_1_2498_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_944 <= bnn_Add_17Sx16S_17S_1_2498_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_945
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_945 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_945 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_945 <= {bnn_N_Mux_64_2_2_1_1636_out1[47], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_945 <= Bline_buffer_48_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_946
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_946 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_946 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_946 <= bnn_N_Mux_2_2_3_1_3337_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_946 <= bnn_N_Mux_2_2_3_1_3337_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_947
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_947 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_947 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_947 <= bnn_N_Mux_2_2_3_1_2140_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_947 <= Bline_buffer_68_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_948
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_948 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_948 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_948 <= bnn_N_Mux_3_2_6_4_1640_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_948 <= Bline_buffer_70_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_949
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_949 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_949 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_949 <= bnn_N_Mux_2_2_3_1_3338_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_949 <= bnn_N_Mux_2_2_3_1_3338_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_950
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_950 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_950 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_950 <= bnn_N_Mux_2_2_3_1_2214_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_950 <= Bline_buffer_90_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_951
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_951 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_951 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_951 <= bnn_N_Muxb_1_2_18_4_236_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_951 <= bnn_N_Muxb_1_2_18_4_236_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_951 <= bnn_Add_17Sx16S_17S_1_2525_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_951 <= bnn_Add_17Sx16S_17S_1_2525_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_952
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_952 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_952 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_952 <= bnn_N_Mux_3_2_6_1_1639_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_952 <= Bline_buffer_49_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_953
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_953 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_953 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_953 <= bnn_N_Mux_2_2_3_1_2196_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_953 <= Bline_buffer_69_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_954
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_954 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_954 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_954 <= {bnn_N_Mux_64_2_2_1_1636_out1[48], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_954 <= Bline_buffer_71_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_955
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_955 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_955 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_955 <= bnn_N_Mux_2_2_3_4_3351_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_955 <= bnn_N_Mux_2_2_3_4_3351_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_956
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_956 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_956 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_956 <= bnn_N_Mux_2_2_3_1_2027_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_956 <= Bline_buffer_91_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_957
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_957 <= 1'b0;
                        end
                     end
                     else begin
                        s_reg_957 <= 1'b0;
                     end
                  end
                  
                  5'd06, 5'd08, 5'd10: begin
                     s_reg_957 <= bnn_N_Muxb_1_2_18_4_237_out1;
                  end
                  
                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        s_reg_957 <= bnn_N_Muxb_1_2_18_4_237_out1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        if (drain1) begin
                        end
                        else begin
                           s_reg_957 <= bnn_Add_17Sx16S_17S_1_2552_out1[16];
                        end
                     end
                     else begin
                        if (bnn_Equal_1Ux1U_1U_1_1_3_out1) begin
                        end
                        else begin
                           s_reg_957 <= bnn_Add_17Sx16S_17S_1_2552_out1[16];
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_958
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_958 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_958 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_958 <= {bnn_N_Mux_64_2_2_1_1636_out1[49], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_958 <= Bline_buffer_72_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_959
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_959 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_959 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_959 <= bnn_N_Mux_2_2_3_1_3365_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_959 <= bnn_N_Mux_2_2_3_1_3365_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_960
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_960 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_960 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_960 <= bnn_N_Mux_2_2_3_1_2044_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_960 <= Bline_buffer_92_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_961
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_961 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_961 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_961 <= {bnn_N_Mux_64_2_2_1_1636_out1[50], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_961 <= Bline_buffer_73_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_962
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_962 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_962 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_962 <= bnn_N_Mux_2_2_3_4_3380_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_962 <= bnn_N_Mux_2_2_3_4_3380_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_963
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_963 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_963 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_963 <= bnn_N_Mux_2_2_3_1_2061_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_963 <= Bline_buffer_93_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_964
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_964 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_964 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_964 <= {bnn_N_Mux_64_2_2_1_1636_out1[51], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_964 <= Bline_buffer_74_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_965
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_965 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_965 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_965 <= bnn_N_Mux_2_2_3_4_3396_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_965 <= bnn_N_Mux_2_2_3_4_3396_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_966
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_966 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_966 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_966 <= bnn_N_Mux_2_2_3_1_2078_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_966 <= Bline_buffer_94_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_967
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_967 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_967 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_967 <= {bnn_N_Mux_64_2_2_1_1636_out1[52], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_967 <= Bline_buffer_75_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_968
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_968 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_968 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_968 <= bnn_N_Mux_2_2_3_4_3412_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_968 <= bnn_N_Mux_2_2_3_4_3412_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_969
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_969 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_969 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_969 <= bnn_N_Mux_2_2_3_1_2095_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_969 <= Bline_buffer_95_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_970
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_970 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_970 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_970 <= {bnn_N_Mux_64_2_2_1_1636_out1[53], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_970 <= Bline_buffer_76_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_971
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_971 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_971 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_971 <= bnn_N_Mux_2_2_3_4_3428_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_971 <= bnn_N_Mux_2_2_3_4_3428_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_972
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_972 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_972 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_972 <= bnn_N_Mux_2_2_3_1_2112_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_972 <= Bline_buffer_96_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_973
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_973 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_973 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_973 <= {bnn_N_Mux_64_2_2_1_1636_out1[54], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_973 <= Bline_buffer_77_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_974
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_974 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_974 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_974 <= bnn_N_Mux_2_2_3_4_3444_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_974 <= bnn_N_Mux_2_2_3_4_3444_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_975
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_975 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_975 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_975 <= bnn_N_Mux_2_2_3_1_2129_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_975 <= Bline_buffer_97_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_976
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_976 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_976 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_976 <= bnn_N_Mux_2_2_3_4_3447_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_976 <= bnn_N_Mux_2_2_3_4_3447_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_977
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_977 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_977 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_977 <= bnn_N_Mux_3_2_6_4_1835_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_977 <= bnn_N_Mux_3_2_6_4_961_out1_slice;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_978
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_978 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_978 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_978 <= {bnn_N_Mux_64_2_2_1_1636_out1[55], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_978 <= Bline_buffer_78_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_979
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_979 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_979 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_979 <= bnn_N_Mux_2_2_3_4_3459_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_979 <= bnn_N_Mux_2_2_3_4_3459_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_980
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_980 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_980 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_980 <= bnn_N_Mux_2_2_3_4_2146_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_980 <= Bline_buffer_98_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_981
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_981 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_981 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_981 <= bnn_N_Mux_3_2_6_1_1642_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_981 <= Bline_buffer_100_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_982
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_982 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_982 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_982 <= bnn_N_Mux_2_2_3_4_3460_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_982 <= bnn_N_Mux_2_2_3_4_3460_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_983
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_983 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_983 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_983 <= bnn_N_Mux_3_2_6_1_1641_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_983 <= Bline_buffer_79_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_984
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_984 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_984 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_984 <= bnn_N_Mux_3_2_6_4_1833_out1_slice;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_984 <= Bline_buffer_99_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_985
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_985 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_985 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_985 <= {bnn_N_Mux_64_2_2_1_1636_out1[56], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_985 <= Bline_buffer_101_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_986
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_986 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_986 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_986 <= bnn_N_Mux_2_2_3_4_3473_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_986 <= bnn_N_Mux_2_2_3_4_3473_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_987
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_987 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_987 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_987 <= {bnn_N_Mux_64_2_2_1_1636_out1[57], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_987 <= Bline_buffer_102_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_988
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_988 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_988 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_988 <= bnn_N_Mux_2_2_3_4_3487_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_988 <= bnn_N_Mux_2_2_3_4_3487_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_989
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_989 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_989 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_989 <= {bnn_N_Mux_64_2_2_1_1636_out1[58], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_989 <= Bline_buffer_103_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_990
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_990 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_990 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_990 <= bnn_N_Mux_2_2_3_4_3502_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_990 <= bnn_N_Mux_2_2_3_4_3502_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_991
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_991 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_991 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_991 <= {bnn_N_Mux_64_2_2_1_1636_out1[59], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_991 <= Bline_buffer_104_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_992
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_992 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_992 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_992 <= bnn_N_Mux_2_2_3_4_3517_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_992 <= bnn_N_Mux_2_2_3_4_3517_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_993
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_993 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_993 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_993 <= {bnn_N_Mux_64_2_2_1_1636_out1[60], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_993 <= Bline_buffer_105_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_994
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_994 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_994 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_994 <= bnn_N_Mux_2_2_3_4_3530_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_994 <= bnn_N_Mux_2_2_3_4_3530_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_995
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_995 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_995 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_995 <= {bnn_N_Mux_64_2_2_1_1636_out1[61], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_995 <= Bline_buffer_106_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_996
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_996 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_996 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_996 <= bnn_N_Mux_2_2_3_4_3539_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_996 <= bnn_N_Mux_2_2_3_4_3539_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_997
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_997 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_997 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_997 <= {bnn_N_Mux_64_2_2_1_1636_out1[62], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_997 <= Bline_buffer_107_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx2i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_998
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_998 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_998 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_998 <= bnn_N_Mux_2_2_3_4_3545_out1;
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           if (cycle2_state) begin
                           end
                           else begin
                              s_reg_998 <= bnn_N_Mux_2_2_3_4_3545_out1;
                           end
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_s_reg_999
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd01: begin
                     if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                        if (32'd0000000000 != s_reg_1005[31:0]) begin
                           s_reg_999 <= 2'd0;
                        end
                     end
                     else begin
                        s_reg_999 <= 2'd0;
                     end
                  end
                  
                  5'd11: begin
                     if (!cycle2_state && !s_reg_1112) begin
                        s_reg_999 <= {bnn_N_Mux_64_2_2_1_1636_out1[63], 1'b1};
                     end
                     else begin
                        if (cycle1_state) begin
                        end
                        else begin
                           s_reg_999 <= Bline_buffer_108_mi61;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: bnn_N_MuxB_160_2_0_4
         always @(xcelreq_data or xcelreq_m_stall_reg_full or xcelreq_m_stall_reg)
          begin :bnn_N_MuxB_160_2_0_4_37
            if (xcelreq_m_stall_reg_full) begin
               bnn_N_MuxB_160_2_0_4_37_out1 = xcelreq_m_stall_reg;
            end
            else begin
               bnn_N_MuxB_160_2_0_4_37_out1 = xcelreq_data;
            end
         end

         assign bnn_Equal_5Ux1U_1U_4_38_in2 = bnn_N_MuxB_160_2_0_4_37_out1[152:148];

         // resource: bnn_Equal_5Ux1U_1U_4  instance: bnn_Equal_5Ux1U_1U_4_38
         assign bnn_Equal_5Ux1U_1U_4_38_out1 = bnn_Equal_5Ux1U_1U_4_38_in2 == 5'd01;

         assign bnn_Equal_7Ux2U_1U_4_39_in2 = {2'b00, bnn_N_MuxB_160_2_0_4_37_out1[152:148]};

         // resource: bnn_Equal_7Ux2U_1U_4  instance: bnn_Equal_7Ux2U_1U_4_39
         assign bnn_Equal_7Ux2U_1U_4_39_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd002;

         // resource: bnn_Equal_7Ux2U_1U_4  instance: bnn_Equal_7Ux2U_1U_4_40
         assign bnn_Equal_7Ux2U_1U_4_40_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd003;

         // resource: bnn_Equal_7Ux3U_1U_4  instance: bnn_Equal_7Ux3U_1U_4_41
         assign bnn_Equal_7Ux3U_1U_4_41_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd004;

         // resource: bnn_Equal_7Ux3U_1U_4  instance: bnn_Equal_7Ux3U_1U_4_42
         assign bnn_Equal_7Ux3U_1U_4_42_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd005;

         // resource: bnn_Equal_7Ux3U_1U_4  instance: bnn_Equal_7Ux3U_1U_4_43
         assign bnn_Equal_7Ux3U_1U_4_43_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd006;

         // resource: mux_5bx2i
         always @(bnn_N_MuxB_160_2_0_4_37_out1[152:148] or bnn_Add_5Sx3S_5S_1_209_out1[3:0] or gs_ctrl4)
          begin :drive_bnn_Equal_5Ux4U_1U_4_44_in2
            if (gs_ctrl4) begin
               bnn_Equal_5Ux4U_1U_4_44_in2 = bnn_N_MuxB_160_2_0_4_37_out1[152:148];
            end
            else begin
               bnn_Equal_5Ux4U_1U_4_44_in2 = {1'b0, bnn_Add_5Sx3S_5S_1_209_out1[3:0]};
            end
         end

         // resource: bnn_Equal_5Ux4U_1U_4  instance: bnn_Equal_5Ux4U_1U_4_44
         assign bnn_Equal_5Ux4U_1U_4_44_out1 = bnn_Equal_5Ux4U_1U_4_44_in2 == 5'd08;

         // resource: bnn_Equal_7Ux3U_1U_4  instance: bnn_Equal_7Ux3U_1U_4_45
         assign bnn_Equal_7Ux3U_1U_4_45_out1 = bnn_Equal_7Ux2U_1U_4_39_in2 == 7'd007;

         assign bnn_Equal_7Ux1U_1U_4_46_in2 = bnn_N_MuxB_160_2_0_4_37_out1[159:153];

         // resource: bnn_Equal_7Ux1U_1U_4  instance: bnn_Equal_7Ux1U_1U_4_46
         assign bnn_Equal_7Ux1U_1U_4_46_out1 = bnn_Equal_7Ux1U_1U_4_46_in2 == 7'd001;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_53
         assign bnn_And_1Sx1U_1U_4_53_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_5Ux1U_1U_4_38_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_54
         assign bnn_And_1Sx1U_1U_4_54_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux2U_1U_4_39_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_55
         assign bnn_And_1Sx1U_1U_4_55_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux2U_1U_4_40_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_56
         assign bnn_And_1Sx1U_1U_4_56_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux3U_1U_4_41_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_57
         assign bnn_And_1Sx1U_1U_4_57_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux3U_1U_4_42_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_58
         assign bnn_And_1Sx1U_1U_4_58_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux3U_1U_4_43_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_59
         assign bnn_And_1Sx1U_1U_4_59_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_5Ux4U_1U_4_44_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_61
         assign bnn_And_1Sx1U_1U_4_61_out1 = bnn_Equal_7Ux1U_1U_4_46_out1 & bnn_Equal_7Ux3U_1U_4_45_out1;

         assign bnn_N_Mux_2_2_3_4_62_in2 = bnn_N_MuxB_160_2_0_4_37_out1[65:64];

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_872 or bnn_And_1Sx1U_1U_4_61_out1 or bnn_N_Mux_2_2_3_4_62_in2)
          begin :bnn_N_Mux_2_2_3_4_62
            if (bnn_And_1Sx1U_1U_4_61_out1) begin
               bnn_N_Mux_2_2_3_4_62_out1 = bnn_N_Mux_2_2_3_4_62_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_4_62_out1 = s_reg_872;
            end
         end

         assign bnn_N_Mux_64_2_2_4_63_in2 = bnn_N_MuxB_160_2_0_4_37_out1[127:64];

         // resource: bnn_N_Mux_64_2_2_4
         always @(s_reg_897 or bnn_And_1Sx1U_1U_4_58_out1 or bnn_N_Mux_64_2_2_4_63_in2)
          begin :bnn_N_Mux_64_2_2_4_63
            if (bnn_And_1Sx1U_1U_4_58_out1) begin
               bnn_N_Mux_64_2_2_4_63_out1 = bnn_N_Mux_64_2_2_4_63_in2;
            end
            else begin
               bnn_N_Mux_64_2_2_4_63_out1 = s_reg_897;
            end
         end

         // resource: bnn_OrReduction_5U_1U_4  instance: bnn_OrReduction_5U_1U_4_64
         assign bnn_OrReduction_5U_1U_4_64_out1 = |bnn_Equal_5Ux1U_1U_4_38_in2;

         // resource: bnn_NotEQ_7Ux1U_1U_4  instance: bnn_NotEQ_7Ux1U_1U_4_65
         assign bnn_NotEQ_7Ux1U_1U_4_65_out1 = bnn_Equal_7Ux1U_1U_4_46_in2 != 7'd001;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_66
         assign bnn_Or_1Sx1U_1S_4_66_out1 = bnn_NotEQ_7Ux1U_1U_4_65_out1 | bnn_OrReduction_5U_1U_4_64_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_67
         assign bnn_And_1Sx1U_1U_4_67_out1 = bnn_Or_1Sx1U_1S_4_66_out1 & s_reg_870;

         assign bnn_N_Muxb_1_2_18_4_68_in2 = bnn_N_MuxB_160_2_0_4_37_out1[64];

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_907 or bnn_And_1Sx1U_1U_4_59_out1 or bnn_N_Muxb_1_2_18_4_68_in2)
          begin :bnn_N_Muxb_1_2_18_4_68
            if (bnn_And_1Sx1U_1U_4_59_out1) begin
               bnn_N_Muxb_1_2_18_4_68_out1 = bnn_N_Muxb_1_2_18_4_68_in2;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_68_out1 = s_reg_907;
            end
         end

         assign bnn_N_Mux_32_2_1_4_69_in2 = bnn_N_MuxB_160_2_0_4_37_out1[95:64];

         // resource: bnn_N_Mux_32_2_1_4
         always @(s_reg_1017 or bnn_And_1Sx1U_1U_4_53_out1 or bnn_N_Mux_32_2_1_4_69_in2)
          begin :bnn_N_Mux_32_2_1_4_69
            if (bnn_And_1Sx1U_1U_4_53_out1) begin
               bnn_N_Mux_32_2_1_4_69_out1 = bnn_N_Mux_32_2_1_4_69_in2;
            end
            else begin
               bnn_N_Mux_32_2_1_4_69_out1 = s_reg_1017;
            end
         end

         // resource: bnn_N_Mux_32_2_1_4
         always @(s_reg_1003 or bnn_And_1Sx1U_1U_4_54_out1 or bnn_N_Mux_32_2_1_4_69_in2)
          begin :bnn_N_Mux_32_2_1_4_70
            if (bnn_And_1Sx1U_1U_4_54_out1) begin
               bnn_N_Mux_32_2_1_4_70_out1 = bnn_N_Mux_32_2_1_4_69_in2;
            end
            else begin
               bnn_N_Mux_32_2_1_4_70_out1 = s_reg_1003;
            end
         end

         // resource: bnn_N_Mux_32_2_1_4
         always @(s_reg_1002 or bnn_And_1Sx1U_1U_4_55_out1 or bnn_N_Mux_32_2_1_4_69_in2)
          begin :bnn_N_Mux_32_2_1_4_71
            if (bnn_And_1Sx1U_1U_4_55_out1) begin
               bnn_N_Mux_32_2_1_4_71_out1 = bnn_N_Mux_32_2_1_4_69_in2;
            end
            else begin
               bnn_N_Mux_32_2_1_4_71_out1 = s_reg_1002;
            end
         end

         // resource: bnn_N_Mux_32_2_1_4
         always @(s_reg_1001 or bnn_And_1Sx1U_1U_4_56_out1 or bnn_N_Mux_32_2_1_4_69_in2)
          begin :bnn_N_Mux_32_2_1_4_72
            if (bnn_And_1Sx1U_1U_4_56_out1) begin
               bnn_N_Mux_32_2_1_4_72_out1 = bnn_N_Mux_32_2_1_4_69_in2;
            end
            else begin
               bnn_N_Mux_32_2_1_4_72_out1 = s_reg_1001;
            end
         end

         // resource: bnn_N_Mux_32_2_1_4
         always @(s_reg_1000 or bnn_And_1Sx1U_1U_4_57_out1 or bnn_N_Mux_32_2_1_4_69_in2)
          begin :bnn_N_Mux_32_2_1_4_73
            if (bnn_And_1Sx1U_1U_4_57_out1) begin
               bnn_N_Mux_32_2_1_4_73_out1 = bnn_N_Mux_32_2_1_4_69_in2;
            end
            else begin
               bnn_N_Mux_32_2_1_4_73_out1 = s_reg_1000;
            end
         end

         // resource: bnn_N_MuxB_64_10_5_4
         always @(bnn_Equal_5Ux1U_1U_4_38_in2 or bnn_N_Mux_2_2_3_4_62_out1 or bnn_N_Mux_64_2_2_4_63_out1 or bnn_N_Muxb_1_2_18_4_68_out1 or bnn_N_Mux_32_2_1_4_69_out1 or bnn_N_Mux_32_2_1_4_70_out1 or bnn_N_Mux_32_2_1_4_71_out1 or bnn_N_Mux_32_2_1_4_72_out1 or bnn_N_Mux_32_2_1_4_73_out1)
          begin :bnn_N_MuxB_64_10_5_4_74
            case (bnn_Equal_5Ux1U_1U_4_38_in2) 

               5'd00: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = 64'd00000000000000000001;
               end
               
               5'd01: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {32'b00000000000000000000000000000000, bnn_N_Mux_32_2_1_4_69_out1};
               end
               
               5'd02: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {32'b00000000000000000000000000000000, bnn_N_Mux_32_2_1_4_70_out1};
               end
               
               5'd03: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {32'b00000000000000000000000000000000, bnn_N_Mux_32_2_1_4_71_out1};
               end
               
               5'd04: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {32'b00000000000000000000000000000000, bnn_N_Mux_32_2_1_4_72_out1};
               end
               
               5'd05: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {32'b00000000000000000000000000000000, bnn_N_Mux_32_2_1_4_73_out1};
               end
               
               5'd06: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = bnn_N_Mux_64_2_2_4_63_out1;
               end
               
               5'd07: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {62'b00000000000000000000000000000000000000000000000000000000000000, bnn_N_Mux_2_2_3_4_62_out1};
               end
               
               5'd08: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = {63'b000000000000000000000000000000000000000000000000000000000000000, bnn_N_Muxb_1_2_18_4_68_out1};
               end
               
               default: begin
                  bnn_N_MuxB_64_10_5_4_74_out1 = 64'd00000000000000000000;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(gs_ctrl198)
          begin :drive_bnn_LeftShift_2Sx2U_5S_4_75_in2
            if (gs_ctrl198) begin
               bnn_LeftShift_2Sx2U_5S_4_75_in2_slice = 1'b0;
            end
            else begin
               bnn_LeftShift_2Sx2U_5S_4_75_in2_slice = 1'b1;
            end
         end

         // resource: bnn_LeftShift_2Sx2U_5S_4  instance: bnn_LeftShift_2Sx2U_5S_4_75
         assign bnn_LeftShift_2Sx2U_5S_4_75_out1 = {{ 4 {bnn_LeftShift_2Sx2U_5S_4_75_in2_slice}}, 1'b1} << s_reg_1004;

         // resource: mux_5bx3i
         always @(bnn_LeftShift_2Sx2U_5S_4_75_out1 or gs_ctrl199)
          begin :drive_bnn_LeftShift_5Sx2U_8S_4_76_in2
            case (gs_ctrl199) 

               2'd1: begin
                  bnn_LeftShift_5Sx2U_8S_4_76_in2 = 5'd31;
               end
               
               2'd2: begin
                  bnn_LeftShift_5Sx2U_8S_4_76_in2 = bnn_LeftShift_2Sx2U_5S_4_75_out1;
               end
               
               default: begin
                  bnn_LeftShift_5Sx2U_8S_4_76_in2 = 5'd08;
               end
               
            endcase

         end

         // resource: bnn_LeftShift_5Sx2U_8S_4  instance: bnn_LeftShift_5Sx2U_8S_4_76
         assign bnn_LeftShift_5Sx2U_8S_4_76_out1 = {{ 3 {bnn_LeftShift_5Sx2U_8S_4_76_in2[4]}}, bnn_LeftShift_5Sx2U_8S_4_76_in2} << s_reg_1004;

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_77
         assign bnn_OrReduction_2U_1U_4_77_out1 = |s_reg_1004;

         // resource: bnn_Equal_2Ux1U_1U_4  instance: bnn_Equal_2Ux1U_1U_4_78
         assign bnn_Equal_2Ux1U_1U_4_78_out1 = s_reg_1004 == 2'd1;

         // resource: bnn_N_Mux_4_2_10_4
         always @(bnn_Equal_2Ux1U_1U_4_78_out1)
          begin :bnn_N_Mux_4_2_10_4_80
            if (bnn_Equal_2Ux1U_1U_4_78_out1) begin
               bnn_N_Mux_4_2_10_4_80_out1_slice = 2'd0;
            end
            else begin
               bnn_N_Mux_4_2_10_4_80_out1_slice = 2'd3;
            end
         end

         // resource: bnn_N_Mux_4_2_11_4
         always @(bnn_OrReduction_2U_1U_4_77_out1 or bnn_N_Mux_4_2_10_4_80_out1_slice)
          begin :bnn_N_Mux_4_2_11_4_83
            if (bnn_OrReduction_2U_1U_4_77_out1) begin
               bnn_N_Mux_4_2_11_4_83_out1 = {bnn_N_Mux_4_2_10_4_80_out1_slice, 2'd3};
            end
            else begin
               bnn_N_Mux_4_2_11_4_83_out1 = 4'd00;
            end
         end

         // resource: bnn_GreaterThan_64Ux10U_1U_4  instance: bnn_GreaterThan_64Ux10U_1U_4_149
         assign bnn_GreaterThan_64Ux10U_1U_4_149_out1 = s_reg_1005 > 64'd00000000000000000512;

         // resource: bnn_GreaterThan_32Ux6U_1U_4  instance: bnn_GreaterThan_32Ux6U_1U_4_179
         assign bnn_GreaterThan_32Ux6U_1U_4_179_out1 = {{ 24 {bnn_LeftShift_5Sx2U_8S_4_76_out1[7]}}, bnn_LeftShift_5Sx2U_8S_4_76_out1} > 32'd0000000032;

         // resource: mux_5bx6i
         always @(s_reg_1027[3:0] or s_reg_1076[4:0] or s_reg_1112 or s_reg_871[3:0] or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_Add_5Sx4S_6S_1_215_out1[4:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or cycle2_state or gs_ctrl205)
          begin :drive_bnn_Add_5Sx4S_6S_1_180_in2
            case (gs_ctrl205) 

               3'd1: begin
                  bnn_Add_5Sx4S_6S_1_180_in2 = {1'b0, s_reg_871[3:0]};
               end
               
               3'd2: begin
                  bnn_Add_5Sx4S_6S_1_180_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
               3'd3: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_180_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_180_in2 = bnn_Add_5Sx4S_6S_1_215_out1[4:0];
                  end
               end
               
               3'd4: begin
                  bnn_Add_5Sx4S_6S_1_180_in2 = {1'b0, s_reg_1027[3:0]};
               end
               
               3'd5: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_180_in2 = bnn_Add_5Sx4S_6S_1_215_out1[4:0];
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_180_in2 = s_reg_1076[4:0];
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_180_in2 = 5'd00;
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_1_1301_out1 or cycle2_state or gs_ctrl206)
          begin :drive_bnn_Add_5Sx4S_6S_1_180_in1
            case (gs_ctrl206) 

               3'd1: begin
                  bnn_Add_5Sx4S_6S_1_180_in1_slice = 3'd0;
               end
               
               3'd2: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_180_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_180_in1_slice = {bnn_N_Mux_2_2_3_1_1301_out1[1], bnn_N_Mux_2_2_3_1_1301_out1};
                  end
               end
               
               3'd3: begin
                  bnn_Add_5Sx4S_6S_1_180_in1_slice = {1'b0, s_reg_1033};
               end
               
               3'd4: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_180_in1_slice = {bnn_N_Mux_2_2_3_1_1301_out1[1], bnn_N_Mux_2_2_3_1_1301_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_180_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_180_in1_slice = 3'd1;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_180
         assign bnn_Add_5Sx4S_6S_1_180_out1 = {bnn_Add_5Sx4S_6S_1_180_in2[4], bnn_Add_5Sx4S_6S_1_180_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_180_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_180_in1_slice};

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_181
         assign bnn_OrReduction_2U_1U_4_181_out1 = |s_reg_1004;

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_189
         assign bnn_OrReduction_2U_1U_4_189_out1 = |s_reg_1004;

         // resource: bnn_LessThan_3Ux3U_1U_4  instance: bnn_LessThan_3Ux3U_1U_4_190
         assign bnn_LessThan_3Ux3U_1U_4_190_out1 = s_reg_1012 < 3'd6;

         // resource: mux_30bx5i
         always @(s_reg_1000[28:0] or s_reg_1003[15:0] or s_reg_1025[1:0] or gs_ctrl210)
          begin :drive_bnn_Mul_30Sx12S_30S_1_191_in2
            case (gs_ctrl210) 

               3'd1: begin
                  bnn_Mul_30Sx12S_30S_1_191_in2 = 30'd0000000000;
               end
               
               3'd2: begin
                  bnn_Mul_30Sx12S_30S_1_191_in2 = {28'b0000000000000000000000000000, s_reg_1025[1:0]};
               end
               
               3'd3: begin
                  bnn_Mul_30Sx12S_30S_1_191_in2 = {1'b0, s_reg_1000[28:0]};
               end
               
               3'd4: begin
                  bnn_Mul_30Sx12S_30S_1_191_in2 = {{ 14 {s_reg_1003[15]}}, s_reg_1003[15:0]};
               end
               
               default: begin
                  bnn_Mul_30Sx12S_30S_1_191_in2 = 30'd0000000009;
               end
               
            endcase

         end

         // resource: mux_12bx4i
         always @(fixed_buffer_0_if_1_dout_wire or s_reg_1012 or s_reg_1019 or gs_ctrl211)
          begin :drive_bnn_Mul_30Sx12S_30S_1_191_in1
            case (gs_ctrl211) 

               2'd1: begin
                  bnn_Mul_30Sx12S_30S_1_191_in1 = 12'd0003;
               end
               
               2'd2: begin
                  bnn_Mul_30Sx12S_30S_1_191_in1 = {2'b00, s_reg_1019};
               end
               
               2'd3: begin
                  bnn_Mul_30Sx12S_30S_1_191_in1 = fixed_buffer_0_if_1_dout_wire;
               end
               
               default: begin
                  bnn_Mul_30Sx12S_30S_1_191_in1 = {9'b000000000, s_reg_1012};
               end
               
            endcase

         end

         // resource: bnn_Mul_30Sx12S_30S_1  instance: bnn_Mul_30Sx12S_30S_1_191
         assign bnn_Mul_30Sx12S_30S_1_191_out1 = bnn_Mul_30Sx12S_30S_1_191_in2*{{ 18 {bnn_Mul_30Sx12S_30S_1_191_in1[11]}}, bnn_Mul_30Sx12S_30S_1_191_in1};

         // resource: mux_10bx2i
         always @(s_reg_1019 or s_reg_1020 or gs_ctrl197)
          begin :drive_bnn_Add_10Ux1U_10U_4_192_in2
            if (gs_ctrl197) begin
               bnn_Add_10Ux1U_10U_4_192_in2 = s_reg_1020;
            end
            else begin
               bnn_Add_10Ux1U_10U_4_192_in2 = s_reg_1019;
            end
         end

         // resource: bnn_Add_10Ux1U_10U_4  instance: bnn_Add_10Ux1U_10U_4_192
         assign bnn_Add_10Ux1U_10U_4_192_out1 = bnn_Add_10Ux1U_10U_4_192_in2 + 10'd0001;

         // resource: mux_6bx6i
         always @(s_reg_1012 or s_reg_1112 or s_reg_871 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_5Sx4S_6S_1_1542_out1[4:0] or cycle2_state or gs_ctrl214)
          begin :drive_bnn_Add_6Sx4S_6S_1_193_in2
            case (gs_ctrl214) 

               3'd1: begin
                  bnn_Add_6Sx4S_6S_1_193_in2 = {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
               3'd2: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_6Sx4S_6S_1_193_in2 = {2'b00, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_6Sx4S_6S_1_193_in2 = {bnn_Add_5Sx4S_6S_1_1542_out1[4], bnn_Add_5Sx4S_6S_1_1542_out1[4:0]};
                  end
               end
               
               3'd3: begin
                  bnn_Add_6Sx4S_6S_1_193_in2 = {2'b00, s_reg_871[3:0]};
               end
               
               3'd4: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_6Sx4S_6S_1_193_in2 = {bnn_Add_5Sx4S_6S_1_1542_out1[4], bnn_Add_5Sx4S_6S_1_1542_out1[4:0]};
                  end
                  else begin
                     bnn_Add_6Sx4S_6S_1_193_in2 = {s_reg_871[4], s_reg_871};
                  end
               end
               
               3'd5: begin
                  bnn_Add_6Sx4S_6S_1_193_in2 = {1'b0, s_reg_871};
               end
               
               default: begin
                  bnn_Add_6Sx4S_6S_1_193_in2 = {3'b000, s_reg_1012};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_4_4057_out1 or cycle2_state or gs_ctrl206)
          begin :drive_bnn_Add_6Sx4S_6S_1_193_in1
            case (gs_ctrl206) 

               3'd1: begin
                  bnn_Add_6Sx4S_6S_1_193_in1_slice = 3'd0;
               end
               
               3'd2: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_6Sx4S_6S_1_193_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_6Sx4S_6S_1_193_in1_slice = {bnn_N_Mux_2_2_3_4_4057_out1[1], bnn_N_Mux_2_2_3_4_4057_out1};
                  end
               end
               
               3'd3: begin
                  bnn_Add_6Sx4S_6S_1_193_in1_slice = {1'b0, s_reg_1033};
               end
               
               3'd4: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_6Sx4S_6S_1_193_in1_slice = {bnn_N_Mux_2_2_3_4_4057_out1[1], bnn_N_Mux_2_2_3_4_4057_out1};
                  end
                  else begin
                     bnn_Add_6Sx4S_6S_1_193_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_6Sx4S_6S_1_193_in1_slice = 3'd1;
               end
               
            endcase

         end

         // resource: bnn_Add_6Sx4S_6S_1  instance: bnn_Add_6Sx4S_6S_1_193
         assign bnn_Add_6Sx4S_6S_1_193_out1 = bnn_Add_6Sx4S_6S_1_193_in2 + {{ 3 {bnn_Add_6Sx4S_6S_1_193_in1_slice[2]}}, bnn_Add_6Sx4S_6S_1_193_in1_slice};

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_194
         assign bnn_OrReduction_2U_1U_4_194_out1 = |s_reg_1004;

         // resource: mux_7bx4i
         always @(s_reg_1025[1:0] or s_reg_1068[4:0] or s_reg_1163[5:0] or gs_ctrl217)
          begin :drive_bnn_Add_7Sx5S_7S_4_195_in2
            case (gs_ctrl217) 

               2'd1: begin
                  bnn_Add_7Sx5S_7S_4_195_in2 = {5'b00000, s_reg_1025[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_7Sx5S_7S_4_195_in2 = {{ 2 {s_reg_1068[4]}}, s_reg_1068[4:0]};
               end
               
               2'd3: begin
                  bnn_Add_7Sx5S_7S_4_195_in2 = {1'b0, s_reg_1163[5:0]};
               end
               
               default: begin
                  bnn_Add_7Sx5S_7S_4_195_in2 = 7'd000;
               end
               
            endcase

         end

         // resource: bnn_Add_7Sx5S_7S_4  instance: bnn_Add_7Sx5S_7S_4_195
         assign bnn_Add_7Sx5S_7S_4_195_out1 = bnn_Add_7Sx5S_7S_4_195_in2 + 7'd001;

         // resource: mux_6bx2i
         always @(s_reg_1021 or s_reg_1133 or gs_ctrl219)
          begin :drive_bnn_Add_6Ux6U_6U_1_206_in2
            if (gs_ctrl219) begin
               bnn_Add_6Ux6U_6U_1_206_in2 = {s_reg_1133[4], s_reg_1133};
            end
            else begin
               bnn_Add_6Ux6U_6U_1_206_in2 = s_reg_1021;
            end
         end

         // resource: mux_5bx3i
         always @(s_reg_1122[1:0] or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_N_Mux_2_2_3_1_3349_out1 or gs_ctrl196)
          begin :drive_bnn_Add_6Ux6U_6U_1_206_in1
            case (gs_ctrl196) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_206_in1_slice = {{ 3 {bnn_N_Mux_2_2_3_1_3349_out1[1]}}, bnn_N_Mux_2_2_3_1_3349_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_206_in1_slice = {{ 3 {s_reg_1122[1]}}, s_reg_1122[1:0]};
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_206_in1_slice = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_206
         assign bnn_Add_6Ux6U_6U_1_206_out1 = bnn_Add_6Ux6U_6U_1_206_in2 + {bnn_Add_6Ux6U_6U_1_206_in1_slice[4], bnn_Add_6Ux6U_6U_1_206_in1_slice};

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_207
         assign bnn_Not_1U_1U_4_207_out1 = !s_reg_1023;

         // resource: mux_2bx2i
         always @(s_reg_1033 or gs_ctrl222)
          begin :drive_bnn_Add_2Ux1U_2U_4_208_in2
            if (gs_ctrl222) begin
               bnn_Add_2Ux1U_2U_4_208_in2 = s_reg_1033;
            end
            else begin
               bnn_Add_2Ux1U_2U_4_208_in2 = 2'd0;
            end
         end

         // resource: bnn_Add_2Ux1U_2U_4  instance: bnn_Add_2Ux1U_2U_4_208
         assign bnn_Add_2Ux1U_2U_4_208_out1 = bnn_Add_2Ux1U_2U_4_208_in2 + 2'd1;

         // resource: mux_5bx4i
         always @(s_reg_1026 or s_reg_1070[3:0] or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or gs_ctrl224)
          begin :drive_bnn_Add_5Sx3S_5S_1_209_in2
            case (gs_ctrl224) 

               2'd1: begin
                  bnn_Add_5Sx3S_5S_1_209_in2 = {1'b0, s_reg_1026};
               end
               
               2'd2: begin
                  bnn_Add_5Sx3S_5S_1_209_in2 = {s_reg_1070[3], s_reg_1070[3:0]};
               end
               
               2'd3: begin
                  bnn_Add_5Sx3S_5S_1_209_in2 = {s_reg_1026[3], s_reg_1026};
               end
               
               default: begin
                  bnn_Add_5Sx3S_5S_1_209_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or gs_ctrl224)
          begin :drive_bnn_Add_5Sx3S_5S_1_209_in1
            case (gs_ctrl224) 

               2'd1: begin
                  bnn_Add_5Sx3S_5S_1_209_in1 = {1'b0, s_reg_1033};
               end
               
               2'd2: begin
                  bnn_Add_5Sx3S_5S_1_209_in1 = 3'd1;
               end
               
               2'd3: begin
                  bnn_Add_5Sx3S_5S_1_209_in1 = {s_reg_1033[1], s_reg_1033};
               end
               
               default: begin
                  bnn_Add_5Sx3S_5S_1_209_in1 = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx3S_5S_1  instance: bnn_Add_5Sx3S_5S_1_209
         assign bnn_Add_5Sx3S_5S_1_209_out1 = bnn_Add_5Sx3S_5S_1_209_in2 + {{ 2 {bnn_Add_5Sx3S_5S_1_209_in1[2]}}, bnn_Add_5Sx3S_5S_1_209_in1};

         // resource: mux_5bx3i
         always @(s_reg_1028 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or gs_ctrl226)
          begin :drive_bnn_Add_5Sx3S_5S_1_211_in2
            case (gs_ctrl226) 

               2'd1: begin
                  bnn_Add_5Sx3S_5S_1_211_in2 = {1'b0, s_reg_1028};
               end
               
               2'd2: begin
                  bnn_Add_5Sx3S_5S_1_211_in2 = {s_reg_1028[3], s_reg_1028};
               end
               
               default: begin
                  bnn_Add_5Sx3S_5S_1_211_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx3i
         always @(s_reg_1033 or bnn_N_Mux_2_2_3_1_3516_out1 or gs_ctrl226)
          begin :drive_bnn_Add_5Sx3S_5S_1_211_in1
            case (gs_ctrl226) 

               2'd1: begin
                  bnn_Add_5Sx3S_5S_1_211_in1 = {1'b0, s_reg_1033};
               end
               
               2'd2: begin
                  bnn_Add_5Sx3S_5S_1_211_in1 = {bnn_N_Mux_2_2_3_1_3516_out1[1], bnn_N_Mux_2_2_3_1_3516_out1};
               end
               
               default: begin
                  bnn_Add_5Sx3S_5S_1_211_in1 = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx3S_5S_1  instance: bnn_Add_5Sx3S_5S_1_211
         assign bnn_Add_5Sx3S_5S_1_211_out1 = bnn_Add_5Sx3S_5S_1_211_in2 + {{ 2 {bnn_Add_5Sx3S_5S_1_211_in1[2]}}, bnn_Add_5Sx3S_5S_1_211_in1};

         // resource: mux_5bx4i
         always @(s_reg_1029[4:0] or s_reg_1112 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_4Sx2S_5S_4_1355_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_212_in2
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_212_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_212_in2 = bnn_Add_4Sx2S_5S_4_1355_out1;
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_212_in2 = {1'b0, s_reg_1029[3:0]};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_212_in2 = bnn_Add_4Sx2S_5S_4_1355_out1;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_212_in2 = s_reg_1029[4:0];
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_212_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_4_4060_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_212_in1
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_212_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_212_in1_slice = {bnn_N_Mux_2_2_3_4_4060_out1[1], bnn_N_Mux_2_2_3_4_4060_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_212_in1_slice = {1'b0, s_reg_1033};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_212_in1_slice = {bnn_N_Mux_2_2_3_4_4060_out1[1], bnn_N_Mux_2_2_3_4_4060_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_212_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_212_in1_slice = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_212
         assign bnn_Add_5Sx4S_6S_1_212_out1 = {bnn_Add_5Sx4S_6S_1_212_in2[4], bnn_Add_5Sx4S_6S_1_212_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_212_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_212_in1_slice};

         // resource: mux_5bx4i
         always @(s_reg_1030 or s_reg_1112 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_4Sx2S_5S_1_1154_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_213_in2
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_213_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_213_in2 = bnn_Add_4Sx2S_5S_1_1154_out1;
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_213_in2 = {1'b0, s_reg_1030[3:0]};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_213_in2 = bnn_Add_4Sx2S_5S_1_1154_out1;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_213_in2 = s_reg_1030;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_213_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_1_1437_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_213_in1
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_213_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_213_in1_slice = {bnn_N_Mux_2_2_3_1_1437_out1[1], bnn_N_Mux_2_2_3_1_1437_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_213_in1_slice = {1'b0, s_reg_1033};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_213_in1_slice = {bnn_N_Mux_2_2_3_1_1437_out1[1], bnn_N_Mux_2_2_3_1_1437_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_213_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_213_in1_slice = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_213
         assign bnn_Add_5Sx4S_6S_1_213_out1 = {bnn_Add_5Sx4S_6S_1_213_in2[4], bnn_Add_5Sx4S_6S_1_213_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_213_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_213_in1_slice};

         // resource: mux_5bx4i
         always @(s_reg_1021[4:0] or s_reg_1036[3:0] or s_reg_1112 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_4Sx2S_5S_1_1261_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_214_in2
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_214_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_214_in2 = bnn_Add_4Sx2S_5S_1_1261_out1;
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_214_in2 = {1'b0, s_reg_1036[3:0]};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_214_in2 = bnn_Add_4Sx2S_5S_1_1261_out1;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_214_in2 = s_reg_1021[4:0];
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_214_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_4_1482_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_214_in1
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_214_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_214_in1_slice = {bnn_N_Mux_2_2_3_4_1482_out1[1], bnn_N_Mux_2_2_3_4_1482_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_214_in1_slice = {1'b0, s_reg_1033};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_214_in1_slice = {bnn_N_Mux_2_2_3_4_1482_out1[1], bnn_N_Mux_2_2_3_4_1482_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_214_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_214_in1_slice = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_214
         assign bnn_Add_5Sx4S_6S_1_214_out1 = {bnn_Add_5Sx4S_6S_1_214_in2[4], bnn_Add_5Sx4S_6S_1_214_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_214_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_214_in1_slice};

         // resource: mux_5bx4i
         always @(s_reg_1031[4:0] or s_reg_1112 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_4Sx2S_5S_1_1269_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_215_in2
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_215_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_215_in2 = bnn_Add_4Sx2S_5S_1_1269_out1;
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_215_in2 = {1'b0, s_reg_1031[3:0]};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_215_in2 = bnn_Add_4Sx2S_5S_1_1269_out1;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_215_in2 = s_reg_1031[4:0];
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_215_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_4_1494_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_215_in1
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_215_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_215_in1_slice = {bnn_N_Mux_2_2_3_4_1494_out1[1], bnn_N_Mux_2_2_3_4_1494_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_215_in1_slice = {1'b0, s_reg_1033};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_215_in1_slice = {bnn_N_Mux_2_2_3_4_1494_out1[1], bnn_N_Mux_2_2_3_4_1494_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_215_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_215_in1_slice = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_215
         assign bnn_Add_5Sx4S_6S_1_215_out1 = {bnn_Add_5Sx4S_6S_1_215_in2[4], bnn_Add_5Sx4S_6S_1_215_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_215_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_215_in1_slice};

         // resource: mux_5bx4i
         always @(s_reg_1035 or s_reg_1112 or bnn_Mul_30Sx12S_30S_1_191_out1[3:0] or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_Add_4Sx2S_5S_1_1280_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_216_in2
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_216_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_216_in2 = bnn_Add_4Sx2S_5S_1_1280_out1;
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_216_in2 = {1'b0, s_reg_1035[3:0]};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_216_in2 = bnn_Add_4Sx2S_5S_1_1280_out1;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_216_in2 = s_reg_1035;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_216_in2 = {1'b0, bnn_Mul_30Sx12S_30S_1_191_out1[3:0]};
               end
               
            endcase

         end

         // resource: mux_3bx4i
         always @(s_reg_1033 or s_reg_1112 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_N_Mux_2_2_3_1_4010_out1 or cycle2_state or gs_ctrl228)
          begin :drive_bnn_Add_5Sx4S_6S_1_216_in1
            case (gs_ctrl228) 

               2'd1: begin
                  if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                     bnn_Add_5Sx4S_6S_1_216_in1_slice = 3'd0;
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_216_in1_slice = {bnn_N_Mux_2_2_3_1_4010_out1[1], bnn_N_Mux_2_2_3_1_4010_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_5Sx4S_6S_1_216_in1_slice = {1'b0, s_reg_1033};
               end
               
               2'd3: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_5Sx4S_6S_1_216_in1_slice = {bnn_N_Mux_2_2_3_1_4010_out1[1], bnn_N_Mux_2_2_3_1_4010_out1};
                  end
                  else begin
                     bnn_Add_5Sx4S_6S_1_216_in1_slice = 3'd1;
                  end
               end
               
               default: begin
                  bnn_Add_5Sx4S_6S_1_216_in1_slice = 3'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_216
         assign bnn_Add_5Sx4S_6S_1_216_out1 = {bnn_Add_5Sx4S_6S_1_216_in2[4], bnn_Add_5Sx4S_6S_1_216_in2} + {{ 3 {bnn_Add_5Sx4S_6S_1_216_in1_slice[2]}}, bnn_Add_5Sx4S_6S_1_216_in1_slice};

         // resource: bnn_Equal_4Ux3U_1U_4  instance: bnn_Equal_4Ux3U_1U_4_219
         assign bnn_Equal_4Ux3U_1U_4_219_out1 = bnn_Add_5Sx4S_6S_1_180_out1[3:0] == 4'd07;

         // resource: bnn_Equal_4Ux3U_1U_4  instance: bnn_Equal_4Ux3U_1U_4_220
         assign bnn_Equal_4Ux3U_1U_4_220_out1 = bnn_Add_5Sx3S_5S_1_211_out1[3:0] == 4'd06;

         // resource: bnn_Equal_4Ux3U_1U_4  instance: bnn_Equal_4Ux3U_1U_4_221
         assign bnn_Equal_4Ux3U_1U_4_221_out1 = bnn_Add_5Sx4S_6S_1_212_out1[3:0] == 4'd05;

         // resource: bnn_Equal_4Ux3U_1U_4  instance: bnn_Equal_4Ux3U_1U_4_222
         assign bnn_Equal_4Ux3U_1U_4_222_out1 = bnn_Add_5Sx4S_6S_1_213_out1[3:0] == 4'd04;

         // resource: bnn_Equal_4Ux2U_1U_4  instance: bnn_Equal_4Ux2U_1U_4_223
         assign bnn_Equal_4Ux2U_1U_4_223_out1 = bnn_Add_5Sx4S_6S_1_214_out1[3:0] == 4'd03;

         // resource: bnn_Equal_4Ux2U_1U_4  instance: bnn_Equal_4Ux2U_1U_4_224
         assign bnn_Equal_4Ux2U_1U_4_224_out1 = bnn_Add_5Sx4S_6S_1_215_out1[3:0] == 4'd02;

         // resource: bnn_Equal_4Ux1U_1U_4  instance: bnn_Equal_4Ux1U_1U_4_225
         assign bnn_Equal_4Ux1U_1U_4_225_out1 = bnn_Add_5Sx4S_6S_1_216_out1[3:0] == 4'd01;

         // resource: bnn_OrReduction_4U_1U_4  instance: bnn_OrReduction_4U_1U_4_226
         assign bnn_OrReduction_4U_1U_4_226_out1 = |bnn_Add_6Sx4S_6S_1_193_out1[3:0];

         // resource: mux_7bx3i
         always @(s_reg_1032 or bnn_Add_6Ux6U_6U_1_206_out1 or gs_ctrl226)
          begin :drive_bnn_Add_7Sx4S_7S_1_227_in2
            case (gs_ctrl226) 

               2'd1: begin
                  bnn_Add_7Sx4S_7S_1_227_in2 = {1'b0, s_reg_1032};
               end
               
               2'd2: begin
                  bnn_Add_7Sx4S_7S_1_227_in2 = {{ 2 {s_reg_1032[4]}}, s_reg_1032[4:0]};
               end
               
               default: begin
                  bnn_Add_7Sx4S_7S_1_227_in2 = {1'b0, bnn_Add_6Ux6U_6U_1_206_out1};
               end
               
            endcase

         end

         // resource: mux_2bx3i
         always @(s_reg_1033 or gs_ctrl226)
          begin :drive_bnn_Add_7Sx4S_7S_1_227_in1
            case (gs_ctrl226) 

               2'd1: begin
                  bnn_Add_7Sx4S_7S_1_227_in1_slice = s_reg_1033;
               end
               
               2'd2: begin
                  bnn_Add_7Sx4S_7S_1_227_in1_slice = 2'd1;
               end
               
               default: begin
                  bnn_Add_7Sx4S_7S_1_227_in1_slice = 2'd0;
               end
               
            endcase

         end

         // resource: bnn_Add_7Sx4S_7S_1  instance: bnn_Add_7Sx4S_7S_1_227
         assign bnn_Add_7Sx4S_7S_1_227_out1 = bnn_Add_7Sx4S_7S_1_227_in2 + {5'd00, bnn_Add_7Sx4S_7S_1_227_in1_slice};

         // resource: mux_64bx3i
         always @(memresp_data[63:0] or s_reg_897 or bnn_N_Mux_64_2_2_1_1636_out1 or gs_ctrl240)
          begin :drive_bnn_RightShift_64Sx8S_1S_1_228_in2
            case (gs_ctrl240) 

               2'd1: begin
                  bnn_RightShift_64Sx8S_1S_1_228_in2 = memresp_data[63:0];
               end
               
               2'd2: begin
                  bnn_RightShift_64Sx8S_1S_1_228_in2 = bnn_N_Mux_64_2_2_1_1636_out1;
               end
               
               default: begin
                  bnn_RightShift_64Sx8S_1S_1_228_in2 = s_reg_897;
               end
               
            endcase

         end

         // resource: mux_8bx2i
         always @(bnn_Add_7Sx4S_7S_1_227_out1[5:0] or gs_ctrl197 or s_reg_1058_stage1_slice[4:0])
          begin :drive_bnn_RightShift_64Sx8S_1S_1_228_in1
            if (gs_ctrl197) begin
               bnn_RightShift_64Sx8S_1S_1_228_in1 = {s_reg_1058_stage1_slice[4:0], 3'd2};
            end
            else begin
               bnn_RightShift_64Sx8S_1S_1_228_in1 = {2'b00, bnn_Add_7Sx4S_7S_1_227_out1[5:0]};
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_228
         assign bnn_RightShift_64Sx8S_1S_1_228_out1 = {{ 64 {bnn_RightShift_64Sx8S_1S_1_228_in2[63]}}, bnn_RightShift_64Sx8S_1S_1_228_in2} >> bnn_RightShift_64Sx8S_1S_1_228_in1[5:0];

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_908 or bnn_Equal_5Ux4U_1U_4_44_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_229
            if (bnn_Equal_5Ux4U_1U_4_44_out1) begin
               bnn_N_Muxb_1_2_18_4_229_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_229_out1 = s_reg_908;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_907 or bnn_Equal_4Ux3U_1U_4_219_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_230
            if (bnn_Equal_4Ux3U_1U_4_219_out1) begin
               bnn_N_Muxb_1_2_18_4_230_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_230_out1 = s_reg_907;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_916 or bnn_Equal_4Ux3U_1U_4_220_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_231
            if (bnn_Equal_4Ux3U_1U_4_220_out1) begin
               bnn_N_Muxb_1_2_18_4_231_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_231_out1 = s_reg_916;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_924 or bnn_Equal_4Ux3U_1U_4_221_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_232
            if (bnn_Equal_4Ux3U_1U_4_221_out1) begin
               bnn_N_Muxb_1_2_18_4_232_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_232_out1 = s_reg_924;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_932 or bnn_Equal_4Ux3U_1U_4_222_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_233
            if (bnn_Equal_4Ux3U_1U_4_222_out1) begin
               bnn_N_Muxb_1_2_18_4_233_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_233_out1 = s_reg_932;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_939 or bnn_Equal_4Ux2U_1U_4_223_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_234
            if (bnn_Equal_4Ux2U_1U_4_223_out1) begin
               bnn_N_Muxb_1_2_18_4_234_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_234_out1 = s_reg_939;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_944 or bnn_Equal_4Ux2U_1U_4_224_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_235
            if (bnn_Equal_4Ux2U_1U_4_224_out1) begin
               bnn_N_Muxb_1_2_18_4_235_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_235_out1 = s_reg_944;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_951 or bnn_Equal_4Ux1U_1U_4_225_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_236
            if (bnn_Equal_4Ux1U_1U_4_225_out1) begin
               bnn_N_Muxb_1_2_18_4_236_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_236_out1 = s_reg_951;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(s_reg_957 or bnn_OrReduction_4U_1U_4_226_out1 or bnn_RightShift_64Sx8S_1S_1_228_out1)
          begin :bnn_N_Muxb_1_2_18_4_237
            if (bnn_OrReduction_4U_1U_4_226_out1) begin
               bnn_N_Muxb_1_2_18_4_237_out1 = s_reg_957;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_237_out1 = bnn_RightShift_64Sx8S_1S_1_228_out1;
            end
         end

         // resource: bnn_LessThan_2Ux2U_1U_4  instance: bnn_LessThan_2Ux2U_1U_4_238
         assign bnn_LessThan_2Ux2U_1U_4_238_out1 = s_reg_1033 < 2'd3;

         // resource: bnn_LessThan_2Ux2U_1U_4  instance: bnn_LessThan_2Ux2U_1U_4_239
         assign bnn_LessThan_2Ux2U_1U_4_239_out1 = s_reg_1025[1:0] < 2'd3;

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_241
         assign bnn_OrReduction_2U_1U_4_241_out1 = |s_reg_1004;

         // resource: bnn_Add_4Sx4S_5S_4  instance: bnn_Add_4Sx4S_5S_4_272
         assign bnn_Add_4Sx4S_5S_4_272_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd04;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1173_out1 or bnn_Mod_3Ux32U_7U_4_4488_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_274_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_274_in2 = {bnn_Add_4Sx2S_5S_1_1173_out1[4], bnn_Add_4Sx2S_5S_1_1173_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_274_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_274_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_274_in2 = bnn_Mod_3Ux32U_7U_4_4488_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_274_in2 = {bnn_Add_4Sx2S_5S_1_1173_out1[4], bnn_Add_4Sx2S_5S_1_1173_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1306_out1 or bnn_LeftShift_9Ux3U_7U_4_4487_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_274_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_274_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1306_out1[1]}}, bnn_N_Mux_2_2_3_1_1306_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_274_in1 = 6'd04;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_274_in1 = 6'd04;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_274_in1 = bnn_LeftShift_9Ux3U_7U_4_4487_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_274_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1306_out1[1]}}, bnn_N_Mux_2_2_3_1_1306_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_274
         assign bnn_Add_6Ux6U_6U_1_274_out1 = bnn_Add_6Ux6U_6U_1_274_in2 + bnn_Add_6Ux6U_6U_1_274_in1;

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_276
         assign bnn_Add_4Sx2S_5S_4_276_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd01;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_278
         assign bnn_GreaterThan_6Sx4S_1U_4_278_out1 = bnn_LeftShift_2Sx2U_5S_4_75_out1[4] ^ bnn_LeftShift_2Sx2U_5S_4_75_out1 > 5'd07;

         // resource: bnn_LessThanEQ_5Sx4S_1U_4  instance: bnn_LessThanEQ_5Sx4S_1U_4_279
         assign bnn_LessThanEQ_5Sx4S_1U_4_279_out1 = bnn_LeftShift_2Sx2U_5S_4_75_out1[4] ^ bnn_LeftShift_2Sx2U_5S_4_75_out1 <= 5'd07;

         // resource: bnn_OrReduction_10U_1U_4  instance: bnn_OrReduction_10U_1U_4_280
         assign bnn_OrReduction_10U_1U_4_280_out1 = |s_reg_1020;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1228_out1 or bnn_Mod_3Ux32U_7U_4_4498_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_282_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_282_in2 = {bnn_Add_4Sx2S_5S_1_1228_out1[4], bnn_Add_4Sx2S_5S_1_1228_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_282_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_282_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_282_in2 = bnn_Mod_3Ux32U_7U_4_4498_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_282_in2 = {bnn_Add_4Sx2S_5S_1_1228_out1[4], bnn_Add_4Sx2S_5S_1_1228_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1450_out1 or bnn_LeftShift_9Ux3U_7U_4_4497_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_282_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_282_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1450_out1[1]}}, bnn_N_Mux_2_2_3_1_1450_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_282_in1 = 6'd01;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_282_in1 = 6'd01;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_282_in1 = bnn_LeftShift_9Ux3U_7U_4_4497_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_282_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1450_out1[1]}}, bnn_N_Mux_2_2_3_1_1450_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_282
         assign bnn_Add_6Ux6U_6U_1_282_out1 = bnn_Add_6Ux6U_6U_1_282_in2 + bnn_Add_6Ux6U_6U_1_282_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_286
         assign bnn_GreaterThan_6Sx4S_1U_4_286_out1 = bnn_Add_4Sx4S_5S_4_272_out1[4] ^ bnn_Add_4Sx4S_5S_4_272_out1 > 5'd07;

         // resource: bnn_LessThanEQ_5Sx4S_1U_4  instance: bnn_LessThanEQ_5Sx4S_1U_4_287
         assign bnn_LessThanEQ_5Sx4S_1U_4_287_out1 = bnn_Add_4Sx4S_5S_4_272_out1[4] ^ bnn_Add_4Sx4S_5S_4_272_out1 <= 5'd07;

         // resource: bnn_Add_4Sx4S_5S_4  instance: bnn_Add_4Sx4S_5S_4_290
         assign bnn_Add_4Sx4S_5S_4_290_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd05;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_294
         assign bnn_GreaterThan_6Sx4S_1U_4_294_out1 = bnn_Add_6Ux6U_6U_1_274_out1[5] ^ bnn_Add_6Ux6U_6U_1_274_out1 > 6'd07;

         // resource: bnn_LessThanEQ_6Sx4S_1U_4  instance: bnn_LessThanEQ_6Sx4S_1U_4_295
         assign bnn_LessThanEQ_6Sx4S_1U_4_295_out1 = bnn_Add_6Ux6U_6U_1_274_out1[5] ^ bnn_Add_6Ux6U_6U_1_274_out1 <= 6'd07;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1245_out1 or bnn_Mod_4Ux32U_7U_4_4508_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_298_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_298_in2 = {bnn_Add_4Sx2S_5S_1_1245_out1[4], bnn_Add_4Sx2S_5S_1_1245_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_298_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_298_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_298_in2 = bnn_Mod_4Ux32U_7U_4_4508_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_298_in2 = {bnn_Add_4Sx2S_5S_1_1245_out1[4], bnn_Add_4Sx2S_5S_1_1245_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1467_out1 or bnn_LeftShift_9Ux3U_7U_4_4507_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_298_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_298_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1467_out1[1]}}, bnn_N_Mux_2_2_3_1_1467_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_298_in1 = 6'd05;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_298_in1 = 6'd05;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_298_in1 = bnn_LeftShift_9Ux3U_7U_4_4507_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_298_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1467_out1[1]}}, bnn_N_Mux_2_2_3_1_1467_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_298
         assign bnn_Add_6Ux6U_6U_1_298_out1 = bnn_Add_6Ux6U_6U_1_298_in2 + bnn_Add_6Ux6U_6U_1_298_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_301
         assign bnn_GreaterThan_6Sx4S_1U_4_301_out1 = bnn_Add_4Sx2S_5S_4_276_out1[4] ^ bnn_Add_4Sx2S_5S_4_276_out1 > 5'd07;

         // resource: bnn_Add_4Sx3S_5S_4  instance: bnn_Add_4Sx3S_5S_4_304
         assign bnn_Add_4Sx3S_5S_4_304_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd03;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_305
         assign bnn_And_1Sx1U_1U_4_305_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_5Sx4S_1U_4_279_out1;

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_307
         assign bnn_Not_1U_1U_4_307_out1 = !bnn_OrReduction_10U_1U_4_280_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_308
         assign bnn_GreaterThan_6Sx4S_1U_4_308_out1 = bnn_Add_6Ux6U_6U_1_282_out1[5] ^ bnn_Add_6Ux6U_6U_1_282_out1 > 6'd07;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1193_out1 or bnn_Mod_3Ux32U_7U_4_4478_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_314_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_314_in2 = {bnn_Add_4Sx2S_5S_1_1193_out1[4], bnn_Add_4Sx2S_5S_1_1193_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_314_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_314_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_314_in2 = bnn_Mod_3Ux32U_7U_4_4478_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_314_in2 = {bnn_Add_4Sx2S_5S_1_1193_out1[4], bnn_Add_4Sx2S_5S_1_1193_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1402_out1 or bnn_LeftShift_9Ux3U_7U_4_4477_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_314_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_314_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1402_out1[1]}}, bnn_N_Mux_2_2_3_1_1402_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_314_in1 = 6'd03;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_314_in1 = 6'd03;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_314_in1 = bnn_LeftShift_9Ux3U_7U_4_4477_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_314_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1402_out1[1]}}, bnn_N_Mux_2_2_3_1_1402_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_314
         assign bnn_Add_6Ux6U_6U_1_314_out1 = bnn_Add_6Ux6U_6U_1_314_in2 + bnn_Add_6Ux6U_6U_1_314_in1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_315
         assign bnn_And_1Sx1U_1U_4_315_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_5Sx4S_1U_4_287_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_318
         assign bnn_GreaterThan_6Sx4S_1U_4_318_out1 = bnn_Add_4Sx4S_5S_4_290_out1[4] ^ bnn_Add_4Sx4S_5S_4_290_out1 > 5'd07;

         // resource: bnn_Add_4Sx4S_5S_4  instance: bnn_Add_4Sx4S_5S_4_323
         assign bnn_Add_4Sx4S_5S_4_323_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd07;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_324
         assign bnn_And_1Sx1U_1U_4_324_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_6Sx4S_1U_4_295_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_327
         assign bnn_GreaterThan_6Sx4S_1U_4_327_out1 = bnn_Add_6Ux6U_6U_1_298_out1[5] ^ bnn_Add_6Ux6U_6U_1_298_out1 > 6'd07;

         // resource: bnn_Sub_32Ux1U_32S_1  instance: bnn_Sub_32Ux1U_32S_1_332
         assign bnn_Sub_32Ux1U_32S_1_332_out1 = s_reg_1000 - 32'd0000000001;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_337
         assign bnn_GreaterThan_6Sx4S_1U_4_337_out1 = bnn_Add_4Sx3S_5S_4_304_out1[4] ^ bnn_Add_4Sx3S_5S_4_304_out1 > 5'd07;

         // resource: bnn_LessThanEQ_5Sx4S_1U_4  instance: bnn_LessThanEQ_5Sx4S_1U_4_338
         assign bnn_LessThanEQ_5Sx4S_1U_4_338_out1 = bnn_Add_4Sx3S_5S_4_304_out1[4] ^ bnn_Add_4Sx3S_5S_4_304_out1 <= 5'd07;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_340
         assign bnn_Or_1Sx1U_1S_4_340_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_278_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_342
         assign bnn_Or_1Sx1U_1S_4_342_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_308_out1;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1125_out1 or bnn_Mod_4Ux32U_7U_4_4518_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_345_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_345_in2 = {bnn_Add_4Sx2S_5S_1_1125_out1[4], bnn_Add_4Sx2S_5S_1_1125_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_345_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_345_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_345_in2 = bnn_Mod_4Ux32U_7U_4_4518_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_345_in2 = {bnn_Add_4Sx2S_5S_1_1125_out1[4], bnn_Add_4Sx2S_5S_1_1125_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1406_out1 or bnn_LeftShift_9Ux3U_7U_4_4517_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_345_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_345_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1406_out1[1]}}, bnn_N_Mux_2_2_3_1_1406_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_345_in1 = 6'd02;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_345_in1 = 6'd02;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_345_in1 = bnn_LeftShift_9Ux3U_7U_4_4517_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_345_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1406_out1[1]}}, bnn_N_Mux_2_2_3_1_1406_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_345
         assign bnn_Add_6Ux6U_6U_1_345_out1 = bnn_Add_6Ux6U_6U_1_345_in2 + bnn_Add_6Ux6U_6U_1_345_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_347
         assign bnn_GreaterThan_6Sx4S_1U_4_347_out1 = bnn_Add_6Ux6U_6U_1_314_out1[5] ^ bnn_Add_6Ux6U_6U_1_314_out1 > 6'd07;

         // resource: bnn_LessThanEQ_6Sx4S_1U_4  instance: bnn_LessThanEQ_6Sx4S_1U_4_348
         assign bnn_LessThanEQ_6Sx4S_1U_4_348_out1 = bnn_Add_6Ux6U_6U_1_314_out1[5] ^ bnn_Add_6Ux6U_6U_1_314_out1 <= 6'd07;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_350
         assign bnn_Or_1Sx1U_1S_4_350_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_286_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_352
         assign bnn_Or_1Sx1U_1S_4_352_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_318_out1;

         // resource: bnn_Add_4Sx4S_5S_4  instance: bnn_Add_4Sx4S_5S_4_355
         assign bnn_Add_4Sx4S_5S_4_355_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd06;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_357
         assign bnn_GreaterThan_6Sx4S_1U_4_357_out1 = bnn_Add_4Sx4S_5S_4_323_out1[4] ^ bnn_Add_4Sx4S_5S_4_323_out1 > 5'd07;

         // resource: bnn_LessThanEQ_5Sx4S_1U_4  instance: bnn_LessThanEQ_5Sx4S_1U_4_358
         assign bnn_LessThanEQ_5Sx4S_1U_4_358_out1 = bnn_Add_4Sx4S_5S_4_323_out1[4] ^ bnn_Add_4Sx4S_5S_4_323_out1 <= 5'd07;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_360
         assign bnn_Or_1Sx1U_1S_4_360_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_294_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_362
         assign bnn_Or_1Sx1U_1S_4_362_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_327_out1;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1137_out1 or bnn_Mod_4Ux32U_7U_4_4528_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_365_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_365_in2 = {bnn_Add_4Sx2S_5S_1_1137_out1[4], bnn_Add_4Sx2S_5S_1_1137_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_365_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_365_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_365_in2 = bnn_Mod_4Ux32U_7U_4_4528_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_365_in2 = {bnn_Add_4Sx2S_5S_1_1137_out1[4], bnn_Add_4Sx2S_5S_1_1137_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_3780_out1 or bnn_LeftShift_9Ux3U_7U_4_4527_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_365_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_365_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3780_out1[1]}}, bnn_N_Mux_2_2_3_1_3780_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_365_in1 = 6'd06;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_365_in1 = 6'd06;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_365_in1 = bnn_LeftShift_9Ux3U_7U_4_4527_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_365_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3780_out1[1]}}, bnn_N_Mux_2_2_3_1_3780_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_365
         assign bnn_Add_6Ux6U_6U_1_365_out1 = bnn_Add_6Ux6U_6U_1_365_in2 + bnn_Add_6Ux6U_6U_1_365_in1;

         // resource: bnn_LessThanEQ_10Ux33U_1U_4  instance: bnn_LessThanEQ_10Ux33U_1U_4_368
         assign bnn_LessThanEQ_10Ux33U_1U_4_368_out1 = {23'b00000000000000000000000, s_reg_1020} <= {bnn_Sub_32Ux1U_32S_1_332_out1[31], bnn_Sub_32Ux1U_32S_1_332_out1};

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_370
         assign bnn_Or_1Sx1U_1S_4_370_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_301_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_374
         assign bnn_And_1Sx1U_1U_4_374_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_5Sx4S_1U_4_338_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_381
         assign bnn_GreaterThan_6Sx4S_1U_4_381_out1 = bnn_Add_6Ux6U_6U_1_345_out1[5] ^ bnn_Add_6Ux6U_6U_1_345_out1 > 6'd07;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_386
         assign bnn_And_1Sx1U_1U_4_386_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_6Sx4S_1U_4_348_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_394
         assign bnn_GreaterThan_6Sx4S_1U_4_394_out1 = bnn_Add_4Sx4S_5S_4_355_out1[4] ^ bnn_Add_4Sx4S_5S_4_355_out1 > 5'd07;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_397
         assign bnn_And_1Sx1U_1U_4_397_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_5Sx4S_1U_4_358_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_405
         assign bnn_GreaterThan_6Sx4S_1U_4_405_out1 = bnn_Add_6Ux6U_6U_1_365_out1[5] ^ bnn_Add_6Ux6U_6U_1_365_out1 > 6'd07;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_4Sx2S_5S_1_1211_out1 or bnn_Mod_3Ux32U_7U_4_4468_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_407_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_407_in2 = {bnn_Add_4Sx2S_5S_1_1211_out1[4], bnn_Add_4Sx2S_5S_1_1211_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_407_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_407_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_407_in2 = bnn_Mod_3Ux32U_7U_4_4468_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_407_in2 = {bnn_Add_4Sx2S_5S_1_1211_out1[4], bnn_Add_4Sx2S_5S_1_1211_out1};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_1_1433_out1 or bnn_LeftShift_9Ux3U_7U_4_4467_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_407_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_407_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1433_out1[1]}}, bnn_N_Mux_2_2_3_1_1433_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_407_in1 = 6'd07;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_407_in1 = 6'd07;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_407_in1 = bnn_LeftShift_9Ux3U_7U_4_4467_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_407_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1433_out1[1]}}, bnn_N_Mux_2_2_3_1_1433_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_407
         assign bnn_Add_6Ux6U_6U_1_407_out1 = bnn_Add_6Ux6U_6U_1_407_in2 + bnn_Add_6Ux6U_6U_1_407_in1;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_6Ux6U_6U_1_345_out1[4:0] or bnn_Mod_4Ux32U_7U_4_4538_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_409_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_409_in2 = {bnn_Add_6Ux6U_6U_1_345_out1[4], bnn_Add_6Ux6U_6U_1_345_out1[4:0]};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_409_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_409_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_409_in2 = bnn_Mod_4Ux32U_7U_4_4538_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_409_in2 = {bnn_Add_6Ux6U_6U_1_345_out1[4], bnn_Add_6Ux6U_6U_1_345_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_4_1292_out1 or bnn_LeftShift_9Ux3U_7U_4_4537_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_409_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_409_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1292_out1[1]}}, bnn_N_Mux_2_2_3_4_1292_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_409_in1 = 6'd60;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_409_in1 = 6'd60;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_409_in1 = bnn_LeftShift_9Ux3U_7U_4_4537_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_409_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1292_out1[1]}}, bnn_N_Mux_2_2_3_4_1292_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_409
         assign bnn_Add_6Ux6U_6U_1_409_out1 = bnn_Add_6Ux6U_6U_1_409_in2 + bnn_Add_6Ux6U_6U_1_409_in1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_427
         assign bnn_Or_1Sx1U_1S_4_427_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_381_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_440
         assign bnn_Or_1Sx1U_1S_4_440_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_394_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_453
         assign bnn_Or_1Sx1U_1S_4_453_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_405_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_454
         assign bnn_GreaterThan_6Sx4S_1U_4_454_out1 = bnn_Add_6Ux6U_6U_1_407_out1[5] ^ bnn_Add_6Ux6U_6U_1_407_out1 > 6'd07;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_6Ux6U_6U_1_365_out1[4:0] or bnn_Mod_4Ux32U_7U_4_4548_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_457_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_457_in2 = {bnn_Add_6Ux6U_6U_1_365_out1[4], bnn_Add_6Ux6U_6U_1_365_out1[4:0]};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_457_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_457_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_457_in2 = bnn_Mod_4Ux32U_7U_4_4548_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_457_in2 = {bnn_Add_6Ux6U_6U_1_365_out1[4], bnn_Add_6Ux6U_6U_1_365_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_4_1471_out1 or bnn_LeftShift_9Ux3U_7U_4_4547_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_457_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_457_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1471_out1[1]}}, bnn_N_Mux_2_2_3_4_1471_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_457_in1 = 6'd61;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_457_in1 = 6'd61;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_457_in1 = bnn_LeftShift_9Ux3U_7U_4_4547_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_457_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1471_out1[1]}}, bnn_N_Mux_2_2_3_4_1471_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_457
         assign bnn_Add_6Ux6U_6U_1_457_out1 = bnn_Add_6Ux6U_6U_1_457_in2 + bnn_Add_6Ux6U_6U_1_457_in1;

         // resource: bnn_Add_4Sx3S_5S_4  instance: bnn_Add_4Sx3S_5S_4_463
         assign bnn_Add_4Sx3S_5S_4_463_out1 = {bnn_LeftShift_5Sx2U_8S_4_76_out1[3], bnn_LeftShift_5Sx2U_8S_4_76_out1[3:0]} + 5'd02;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_465
         assign bnn_Or_1Sx1U_1S_4_465_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_337_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_476
         assign bnn_Or_1Sx1U_1S_4_476_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_347_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_487
         assign bnn_Or_1Sx1U_1S_4_487_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_357_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_498
         assign bnn_Or_1Sx1U_1S_4_498_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_454_out1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_503
         assign bnn_GreaterThan_6Sx4S_1U_4_503_out1 = bnn_Add_4Sx3S_5S_4_463_out1[4] ^ bnn_Add_4Sx3S_5S_4_463_out1 > 5'd07;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_550
         assign bnn_Or_1Sx1U_1S_4_550_out1 = bnn_Not_1U_1U_4_307_out1 | bnn_GreaterThan_6Sx4S_1U_4_503_out1;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_5Sx4S_6S_1_213_out1[4:0] or bnn_Mod_4Ux32U_7U_4_4558_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_699_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_699_in2 = {bnn_Add_5Sx4S_6S_1_213_out1[4], bnn_Add_5Sx4S_6S_1_213_out1[4:0]};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_699_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_699_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_699_in2 = bnn_Mod_4Ux32U_7U_4_4558_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_699_in2 = {bnn_Add_5Sx4S_6S_1_213_out1[4], bnn_Add_5Sx4S_6S_1_213_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_4_3827_out1 or bnn_LeftShift_9Ux3U_7U_4_4557_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_699_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_699_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3827_out1[1]}}, bnn_N_Mux_2_2_3_4_3827_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_699_in1 = 6'd62;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_699_in1 = 6'd62;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_699_in1 = bnn_LeftShift_9Ux3U_7U_4_4557_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_699_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3827_out1[1]}}, bnn_N_Mux_2_2_3_4_3827_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_699
         assign bnn_Add_6Ux6U_6U_1_699_out1 = bnn_Add_6Ux6U_6U_1_699_in2 + bnn_Add_6Ux6U_6U_1_699_in1;

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_700
         assign bnn_OrReduction_2U_1U_4_700_out1 = |s_reg_1004;

         // resource: bnn_NotEQ_2Ux1U_1U_4  instance: bnn_NotEQ_2Ux1U_1U_4_701
         assign bnn_NotEQ_2Ux1U_1U_4_701_out1 = s_reg_1004 != 2'd1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_737
         assign bnn_And_1Sx1U_1U_4_737_out1 = bnn_NotEQ_2Ux1U_1U_4_701_out1 & bnn_OrReduction_2U_1U_4_700_out1;

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_LeftShift_2Sx2U_5S_4_75_out1 or bnn_Add_5Sx4S_6S_1_214_out1[4:0] or bnn_Mod_4Ux32U_7U_4_4568_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_887_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_887_in2 = {bnn_Add_5Sx4S_6S_1_214_out1[4], bnn_Add_5Sx4S_6S_1_214_out1[4:0]};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_887_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_887_in2 = {bnn_LeftShift_2Sx2U_5S_4_75_out1[4], bnn_LeftShift_2Sx2U_5S_4_75_out1};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_887_in2 = bnn_Mod_4Ux32U_7U_4_4568_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_887_in2 = {bnn_Add_5Sx4S_6S_1_214_out1[4], bnn_Add_5Sx4S_6S_1_214_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(drain2 or s_reg_1112 or bnn_N_Mux_2_2_3_4_1491_out1 or bnn_LeftShift_9Ux3U_7U_4_4567_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_887_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     if (drain2) begin
                        bnn_Add_6Ux6U_6U_1_887_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1491_out1[1]}}, bnn_N_Mux_2_2_3_4_1491_out1};
                     end
                     else begin
                        bnn_Add_6Ux6U_6U_1_887_in1 = 6'd63;
                     end
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_887_in1 = 6'd63;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_887_in1 = bnn_LeftShift_9Ux3U_7U_4_4567_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_887_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1491_out1[1]}}, bnn_N_Mux_2_2_3_4_1491_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_887
         assign bnn_Add_6Ux6U_6U_1_887_out1 = bnn_Add_6Ux6U_6U_1_887_in2 + bnn_Add_6Ux6U_6U_1_887_in1;

         // resource: bnn_LessThanEQ_6Sx4S_1U_4  instance: bnn_LessThanEQ_6Sx4S_1U_4_950
         assign bnn_LessThanEQ_6Sx4S_1U_4_950_out1 = bnn_Add_6Ux6U_6U_1_407_out1[5] ^ bnn_Add_6Ux6U_6U_1_407_out1 <= 6'd07;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_952
         assign bnn_And_1Sx1U_1U_4_952_out1 = bnn_OrReduction_10U_1U_4_280_out1 & bnn_LessThanEQ_6Sx4S_1U_4_950_out1;

         // resource: mux_32bx4i
         always @(s_reg_1010 or s_reg_1017 or bnn_Mul_30Sx12S_30S_1_191_out1[28:0] or gs_ctrl264)
          begin :drive_bnn_Add_32Ux10U_32U_1_954_in2
            case (gs_ctrl264) 

               2'd1: begin
                  bnn_Add_32Ux10U_32U_1_954_in2 = s_reg_1017;
               end
               
               2'd2: begin
                  bnn_Add_32Ux10U_32U_1_954_in2 = {3'b000, s_reg_1017[28:0]};
               end
               
               2'd3: begin
                  bnn_Add_32Ux10U_32U_1_954_in2 = s_reg_1010;
               end
               
               default: begin
                  bnn_Add_32Ux10U_32U_1_954_in2 = {3'b000, bnn_Mul_30Sx12S_30S_1_191_out1[28:0]};
               end
               
            endcase

         end

         // resource: mux_10bx4i
         always @(s_reg_1020 or s_reg_1024 or s_reg_871 or bnn_Equal_2Ux2U_1U_4_4460_out1 or gs_ctrl264)
          begin :drive_bnn_Add_32Ux10U_32U_1_954_in1
            case (gs_ctrl264) 

               2'd1: begin
                  bnn_Add_32Ux10U_32U_1_954_in1 = {{6'b000000, s_reg_1024}, 3'd0};
               end
               
               2'd2: begin
                  bnn_Add_32Ux10U_32U_1_954_in1 = {9'b000000000, bnn_Equal_2Ux2U_1U_4_4460_out1};
               end
               
               2'd3: begin
                  bnn_Add_32Ux10U_32U_1_954_in1 = {{2'b00, s_reg_871}, 3'd0};
               end
               
               default: begin
                  bnn_Add_32Ux10U_32U_1_954_in1 = s_reg_1020;
               end
               
            endcase

         end

         // resource: bnn_Add_32Ux10U_32U_1  instance: bnn_Add_32Ux10U_32U_1_954
         assign bnn_Add_32Ux10U_32U_1_954_out1 = bnn_Add_32Ux10U_32U_1_954_in2 + {22'b0000000000000000000000, bnn_Add_32Ux10U_32U_1_954_in1};

         // resource: mux_32bx3i
         always @(drain1 or s_reg_1011 or s_reg_1017[28:0] or bnn_Add_32Ux10U_32U_1_954_out1[28:0] or s_reg_1044_stage2 or cycle3_state or gs_ctrl266)
          begin :drive_bnn_Add_32Ux32U_32U_1_955_in2
            case (gs_ctrl266) 

               2'd1: begin
                  bnn_Add_32Ux32U_32U_1_955_in2 = s_reg_1011;
               end
               
               2'd2: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        bnn_Add_32Ux32U_32U_1_955_in2 = s_reg_1011;
                     end
                     else begin
                        bnn_Add_32Ux32U_32U_1_955_in2 = {s_reg_1017[28:0], 3'd0};
                     end
                  end
                  else begin
                     bnn_Add_32Ux32U_32U_1_955_in2 = {s_reg_1017[28:0], 3'd0};
                  end
               end
               
               default: begin
                  bnn_Add_32Ux32U_32U_1_955_in2 = {bnn_Add_32Ux10U_32U_1_954_out1[28:0], 3'd0};
               end
               
            endcase

         end

         // resource: mux_32bx5i
         always @(drain1 or s_reg_1009 or s_reg_1010 or s_reg_871[3:0] or s_reg_886[3:0] or bnn_Add_7Sx5S_7S_4_195_out1 or s_reg_1044_stage2 or cycle3_state or gs_ctrl267)
          begin :drive_bnn_Add_32Ux32U_32U_1_955_in1
            case (gs_ctrl267) 

               2'd1: begin
                  bnn_Add_32Ux32U_32U_1_955_in1 = 32'd0000000000;
               end
               
               2'd2: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     if (drain1) begin
                        bnn_Add_32Ux32U_32U_1_955_in1 = 32'd0000000000;
                     end
                     else begin
                        bnn_Add_32Ux32U_32U_1_955_in1 = s_reg_1010;
                     end
                  end
                  else begin
                     bnn_Add_32Ux32U_32U_1_955_in1 = s_reg_1010;
                  end
               end
               
               2'd3: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     bnn_Add_32Ux32U_32U_1_955_in1 = {{19'b0000000000000000000, s_reg_886[3:0]}, 9'd000};
                  end
                  else begin
                     bnn_Add_32Ux32U_32U_1_955_in1 = {{{19'b0000000000000000000, s_reg_871[3:0]}, bnn_Add_7Sx5S_7S_4_195_out1[5:0]}, 3'd0};
                  end
               end
               
               default: begin
                  bnn_Add_32Ux32U_32U_1_955_in1 = s_reg_1009;
               end
               
            endcase

         end

         // resource: bnn_Add_32Ux32U_32U_1  instance: bnn_Add_32Ux32U_32U_1_955
         assign bnn_Add_32Ux32U_32U_1_955_out1 = bnn_Add_32Ux32U_32U_1_955_in2 + bnn_Add_32Ux32U_32U_1_955_in1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_956
         assign bnn_And_1Sx1U_1U_4_956_out1 = s_reg_1071 & s_reg_1064;

         assign bnn_N_Mux_3_2_6_4_957_ctrl1 = s_reg_1068[5];

         // resource: bnn_N_Mux_3_2_6_4
         always @(Bline_buffer_20_mi61 or bnn_N_Mux_3_2_6_4_957_ctrl1)
          begin :bnn_N_Mux_3_2_6_4_957
            if (bnn_N_Mux_3_2_6_4_957_ctrl1) begin
               bnn_N_Mux_3_2_6_4_957_out1_slice = Bline_buffer_20_mi61;
            end
            else begin
               bnn_N_Mux_3_2_6_4_957_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_7_4
         always @(Bline_buffer_0_mi61 or Bline_buffer_30_mi61 or s_reg_1004 or bnn_N_Mux_3_2_6_4_957_out1_slice)
          begin :bnn_N_Mux_2_4_7_4_958
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_7_4_958_out1 = bnn_N_Mux_3_2_6_4_957_out1_slice;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_7_4_958_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_7_4_958_out1 = Bline_buffer_0_mi61;
               end
               
               default: begin
                  bnn_N_Mux_2_4_7_4_958_out1 = Bline_buffer_30_mi61;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_956_out1 or bnn_N_Mux_2_4_7_4_958_out1)
          begin :bnn_N_Mux_3_2_6_4_959
            if (bnn_And_1Sx1U_1U_4_956_out1) begin
               bnn_N_Mux_3_2_6_4_959_out1_slice = bnn_N_Mux_2_4_7_4_958_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_959_out1_slice = 2'd0;
            end
         end

         // resource: mux_2bx3i
         always @(s_reg_1112 or s_reg_955 or bnn_N_Mux_2_2_3_4_3351_out1 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_959_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_960_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_960_in1 = bnn_N_Mux_2_2_3_4_3351_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_960_in1 = bnn_N_Mux_3_2_6_4_959_out1_slice;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_960_in1 = s_reg_955;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_960
         assign bnn_Minus_2S_2S_4_960_out1 = -bnn_Minus_2S_2S_4_960_in1;

         assign bnn_N_Mux_3_2_6_4_961_ctrl1 = s_reg_1093[5];

         // resource: bnn_N_Mux_3_2_6_4
         always @(Bline_buffer_119_mi61 or bnn_N_Mux_3_2_6_4_961_ctrl1)
          begin :bnn_N_Mux_3_2_6_4_961
            if (bnn_N_Mux_3_2_6_4_961_ctrl1) begin
               bnn_N_Mux_3_2_6_4_961_out1_slice = Bline_buffer_119_mi61;
            end
            else begin
               bnn_N_Mux_3_2_6_4_961_out1_slice = 2'd0;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_1_mi61 or s_reg_1112 or s_reg_874[1:0] or bnn_N_Mux_2_2_3_1_1831_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_962_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_962_in1 = bnn_N_Mux_2_2_3_1_1831_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_962_in1 = Bline_buffer_1_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_962_in1 = s_reg_874[1:0];
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_962
         assign bnn_Minus_2S_2S_1_962_out1 = -bnn_Minus_2S_2S_1_962_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_0_mi61 or s_reg_1112 or s_reg_887 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_963_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_963_in1 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_963_in1 = Bline_buffer_0_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_963_in1 = s_reg_887;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_963
         assign bnn_Minus_2S_2S_4_963_out1 = -bnn_Minus_2S_2S_4_963_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_2_mi61 or s_reg_1112 or s_reg_875 or s_reg_972 or bnn_N_Mux_2_2_3_1_1846_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_964_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_964_in1 = bnn_N_Mux_2_2_3_1_1846_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_964_in1 = Bline_buffer_2_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_964_in1 = s_reg_972;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_964_in1 = s_reg_875;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_964
         assign bnn_Minus_2S_2S_1_964_out1 = -bnn_Minus_2S_2S_1_964_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_1_mi61 or s_reg_1112 or s_reg_874[1:0] or s_reg_969 or bnn_N_Mux_2_2_3_1_1831_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_965_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_965_in1 = bnn_N_Mux_2_2_3_1_1831_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_965_in1 = Bline_buffer_1_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_965_in1 = s_reg_969;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_965_in1 = s_reg_874[1:0];
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_965
         assign bnn_Minus_2S_2S_1_965_out1 = -bnn_Minus_2S_2S_1_965_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_1_mi61 or s_reg_1112 or s_reg_874[1:0] or bnn_N_Mux_2_2_3_1_1831_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_966_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_966_in3 = bnn_N_Mux_2_2_3_1_1831_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_966_in3 = Bline_buffer_1_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_966_in3 = s_reg_874[1:0];
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_Minus_2S_2S_1_962_out1 or bnn_N_Mux_2_2_3_4_966_in3)
          begin :bnn_N_Mux_2_2_3_4_966
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_966_out1 = bnn_Minus_2S_2S_1_962_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_966_out1 = bnn_N_Mux_2_2_3_4_966_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_0_mi61 or s_reg_1112 or s_reg_887 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_967_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_967_in3 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_967_in3 = Bline_buffer_0_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_967_in3 = s_reg_887;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_Minus_2S_2S_4_963_out1 or bnn_N_Mux_2_2_3_4_967_in3)
          begin :bnn_N_Mux_2_2_3_4_967
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_967_out1 = bnn_Minus_2S_2S_4_963_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_967_out1 = bnn_N_Mux_2_2_3_4_967_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_2_mi61 or s_reg_1112 or s_reg_875 or s_reg_996 or bnn_N_Mux_2_2_3_1_1846_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_968_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_968_in1 = bnn_N_Mux_2_2_3_1_1846_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_968_in1 = Bline_buffer_2_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_968_in1 = s_reg_996;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_968_in1 = s_reg_875;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_968
         assign bnn_Minus_2S_2S_1_968_out1 = -bnn_Minus_2S_2S_1_968_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_2_mi61 or s_reg_1112 or s_reg_875 or s_reg_972 or bnn_N_Mux_2_2_3_1_1846_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_969_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_969_in3 = bnn_N_Mux_2_2_3_1_1846_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_969_in3 = Bline_buffer_2_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_969_in3 = s_reg_972;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_969_in3 = s_reg_875;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_964_out1 or bnn_N_Mux_2_2_3_1_969_in3)
          begin :bnn_N_Mux_2_2_3_1_969
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_969_out1 = bnn_Minus_2S_2S_1_964_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_969_out1 = bnn_N_Mux_2_2_3_1_969_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_1_mi61 or s_reg_1112 or s_reg_874[1:0] or s_reg_969 or bnn_N_Mux_2_2_3_1_1831_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_970_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_970_in3 = bnn_N_Mux_2_2_3_1_1831_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_970_in3 = Bline_buffer_1_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_970_in3 = s_reg_969;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_970_in3 = s_reg_874[1:0];
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_965_out1 or bnn_N_Mux_2_2_3_1_970_in3)
          begin :bnn_N_Mux_2_2_3_1_970
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_970_out1 = bnn_Minus_2S_2S_1_965_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_970_out1 = bnn_N_Mux_2_2_3_1_970_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_3_mi61 or s_reg_1112 or s_reg_881 or s_reg_975 or bnn_N_Mux_2_2_3_1_1857_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_971_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_971_in1 = bnn_N_Mux_2_2_3_1_1857_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_971_in1 = Bline_buffer_3_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_971_in1 = s_reg_975;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_971_in1 = s_reg_881;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_971
         assign bnn_Minus_2S_2S_1_971_out1 = -bnn_Minus_2S_2S_1_971_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_972
         assign bnn_Minus_2S_2S_1_972_out1 = -bnn_Minus_2S_2S_1_971_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_973
         assign bnn_Minus_2S_2S_1_973_out1 = -bnn_Minus_2S_2S_1_964_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_11_mi61 or s_reg_1112 or s_reg_876 or bnn_N_Mux_64_2_2_1_1636_out1[32] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_974_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_974_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_974_in1 = Bline_buffer_11_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_974_in1 = s_reg_876;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_974
         assign bnn_Minus_2S_2S_4_974_out1 = -bnn_Minus_2S_2S_4_974_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_975
         assign bnn_Add_2Sx2S_3S_1_975_out1 = {bnn_N_Mux_2_2_3_4_967_out1[1], bnn_N_Mux_2_2_3_4_967_out1} + {bnn_N_Mux_2_2_3_4_966_out1[1], bnn_N_Mux_2_2_3_4_966_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_2_mi61 or s_reg_1112 or s_reg_875 or s_reg_996 or bnn_N_Mux_2_2_3_1_1846_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_976_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_976_in3 = bnn_N_Mux_2_2_3_1_1846_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_976_in3 = Bline_buffer_2_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_976_in3 = s_reg_996;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_976_in3 = s_reg_875;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_916 or s_reg_957 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_976_ctrl1
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_976_ctrl1 = s_reg_957;
            end
            else begin
               bnn_N_Mux_2_2_3_1_976_ctrl1 = s_reg_916;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_968_out1 or bnn_N_Mux_2_2_3_1_976_in3 or bnn_N_Mux_2_2_3_1_976_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_976
            if (bnn_N_Mux_2_2_3_1_976_ctrl1) begin
               bnn_N_Mux_2_2_3_1_976_out1 = bnn_Minus_2S_2S_1_968_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_976_out1 = bnn_N_Mux_2_2_3_1_976_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_11_mi61 or s_reg_1112 or s_reg_876 or s_reg_993 or bnn_N_Mux_64_2_2_1_1636_out1[32] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_977_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_977_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_977_in1 = Bline_buffer_11_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_977_in1 = s_reg_993;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_977_in1 = s_reg_876;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_977
         assign bnn_Minus_2S_2S_1_977_out1 = -bnn_Minus_2S_2S_1_977_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_978
         assign bnn_Add_2Sx2S_3S_1_978_out1 = {bnn_N_Mux_2_2_3_1_970_out1[1], bnn_N_Mux_2_2_3_1_970_out1} + {bnn_N_Mux_2_2_3_1_969_out1[1], bnn_N_Mux_2_2_3_1_969_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_3_mi61 or s_reg_1112 or s_reg_881 or s_reg_975 or bnn_N_Mux_2_2_3_1_1857_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_979_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_979_in3 = bnn_N_Mux_2_2_3_1_1857_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_979_in3 = Bline_buffer_3_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_979_in3 = s_reg_975;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_979_in3 = s_reg_881;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_971_out1 or bnn_N_Mux_2_2_3_1_979_in3)
          begin :bnn_N_Mux_2_2_3_1_979
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_979_out1 = bnn_Minus_2S_2S_1_971_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_979_out1 = bnn_N_Mux_2_2_3_1_979_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_972_out1 or bnn_N_Mux_2_2_3_1_979_in3)
          begin :bnn_N_Mux_2_2_3_1_980
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_980_out1 = bnn_Minus_2S_2S_1_972_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_980_out1 = bnn_N_Mux_2_2_3_1_979_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_969_in3 or bnn_Minus_2S_2S_1_973_out1)
          begin :bnn_N_Mux_2_2_3_1_981
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_981_out1 = bnn_Minus_2S_2S_1_973_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_981_out1 = bnn_N_Mux_2_2_3_1_969_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_4_mi61 or s_reg_1112 or s_reg_888 or s_reg_980 or bnn_N_Mux_2_2_3_1_1868_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_982_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_982_in1 = bnn_N_Mux_2_2_3_1_1868_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_982_in1 = Bline_buffer_4_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_982_in1 = s_reg_980;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_982_in1 = s_reg_888;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_982
         assign bnn_Minus_2S_2S_1_982_out1 = -bnn_Minus_2S_2S_1_982_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_983
         assign bnn_Minus_2S_2S_1_983_out1 = -bnn_Minus_2S_2S_1_982_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_984
         assign bnn_Minus_2S_2S_1_984_out1 = -bnn_Minus_2S_2S_1_971_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_12_mi61 or s_reg_1112 or s_reg_877 or bnn_N_Mux_64_2_2_1_1636_out1[33] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_985_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_985_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_985_in1 = Bline_buffer_12_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_985_in1 = s_reg_877;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_985
         assign bnn_Minus_2S_2S_4_985_out1 = -bnn_Minus_2S_2S_4_985_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_11_mi61 or s_reg_1112 or s_reg_876 or bnn_N_Mux_64_2_2_1_1636_out1[32] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_986_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_986_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_986_in3 = Bline_buffer_11_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_986_in3 = s_reg_876;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_974_out1 or bnn_N_Mux_2_2_3_4_986_in3)
          begin :bnn_N_Mux_2_2_3_4_986
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_986_out1 = bnn_Minus_2S_2S_4_974_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_986_out1 = bnn_N_Mux_2_2_3_4_986_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_987
         assign bnn_Add_3Sx3S_4S_4_987_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_976_out1[1]}}, bnn_N_Mux_2_2_3_1_976_out1} + {bnn_Add_2Sx2S_3S_1_975_out1[2], bnn_Add_2Sx2S_3S_1_975_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_12_mi61 or s_reg_1112 or s_reg_877 or s_reg_995 or bnn_N_Mux_64_2_2_1_1636_out1[33] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_988_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_988_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_988_in1 = Bline_buffer_12_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_988_in1 = s_reg_995;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_988_in1 = s_reg_877;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_988
         assign bnn_Minus_2S_2S_1_988_out1 = -bnn_Minus_2S_2S_1_988_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_11_mi61 or s_reg_1112 or s_reg_876 or s_reg_993 or bnn_N_Mux_64_2_2_1_1636_out1[32] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_989_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_989_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_989_in3 = Bline_buffer_11_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_989_in3 = s_reg_993;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_989_in3 = s_reg_876;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_977_out1 or bnn_N_Mux_2_2_3_1_989_in3)
          begin :bnn_N_Mux_2_2_3_1_989
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_989_out1 = bnn_Minus_2S_2S_1_977_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_989_out1 = bnn_N_Mux_2_2_3_1_989_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_990
         assign bnn_Add_3Sx3S_4S_1_990_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_979_out1[1]}}, bnn_N_Mux_2_2_3_1_979_out1} + {bnn_Add_2Sx2S_3S_1_978_out1[2], bnn_Add_2Sx2S_3S_1_978_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_991
         assign bnn_Minus_2S_2S_1_991_out1 = -bnn_Minus_2S_2S_1_988_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_992
         assign bnn_Add_2Sx2S_3S_1_992_out1 = {bnn_N_Mux_2_2_3_1_981_out1[1], bnn_N_Mux_2_2_3_1_981_out1} + {bnn_N_Mux_2_2_3_1_980_out1[1], bnn_N_Mux_2_2_3_1_980_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_4_mi61 or s_reg_1112 or s_reg_888 or s_reg_980 or bnn_N_Mux_2_2_3_1_1868_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_993_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_993_in3 = bnn_N_Mux_2_2_3_1_1868_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_993_in3 = Bline_buffer_4_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_993_in3 = s_reg_980;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_993_in3 = s_reg_888;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_982_out1 or bnn_N_Mux_2_2_3_1_993_in3)
          begin :bnn_N_Mux_2_2_3_1_993
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_993_out1 = bnn_Minus_2S_2S_1_982_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_993_out1 = bnn_N_Mux_2_2_3_1_993_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_983_out1 or bnn_N_Mux_2_2_3_1_993_in3)
          begin :bnn_N_Mux_2_2_3_1_994
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_994_out1 = bnn_Minus_2S_2S_1_983_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_994_out1 = bnn_N_Mux_2_2_3_1_993_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_979_in3 or bnn_Minus_2S_2S_1_984_out1)
          begin :bnn_N_Mux_2_2_3_1_995
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_995_out1 = bnn_Minus_2S_2S_1_984_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_995_out1 = bnn_N_Mux_2_2_3_1_979_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_5_mi61 or s_reg_1112 or s_reg_898 or s_reg_984 or bnn_N_Mux_2_2_3_1_1879_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_996_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_996_in1 = bnn_N_Mux_2_2_3_1_1879_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_996_in1 = Bline_buffer_5_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_996_in1 = s_reg_984;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_996_in1 = s_reg_898;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_996
         assign bnn_Minus_2S_2S_1_996_out1 = -bnn_Minus_2S_2S_1_996_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_5_mi61 or s_reg_1112 or s_reg_898 or bnn_N_Mux_2_2_3_1_1879_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_997_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_997_in1 = bnn_N_Mux_2_2_3_1_1879_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_997_in1 = Bline_buffer_5_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_997_in1 = s_reg_898;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_997
         assign bnn_Minus_2S_2S_1_997_out1 = -bnn_Minus_2S_2S_1_997_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_4_mi61 or s_reg_1112 or s_reg_888 or bnn_N_Mux_2_2_3_1_1868_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_998_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_998_in1 = bnn_N_Mux_2_2_3_1_1868_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_998_in1 = Bline_buffer_4_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_998_in1 = s_reg_888;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_998
         assign bnn_Minus_2S_2S_1_998_out1 = -bnn_Minus_2S_2S_1_998_in1;

         // resource: mux_2bx3i
         always @(s_reg_1112 or s_reg_959 or bnn_N_Mux_2_2_3_1_3365_out1 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_957_out1_slice)
          begin :drive_bnn_Minus_2S_2S_1_999_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_999_in1 = bnn_N_Mux_2_2_3_1_3365_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_999_in1 = bnn_N_Mux_3_2_6_4_957_out1_slice;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_999_in1 = s_reg_959;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_999
         assign bnn_Minus_2S_2S_1_999_out1 = -bnn_Minus_2S_2S_1_999_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_12_mi61 or s_reg_1112 or s_reg_877 or bnn_N_Mux_64_2_2_1_1636_out1[33] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1000_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1000_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1000_in3 = Bline_buffer_12_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1000_in3 = s_reg_877;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_985_out1 or bnn_N_Mux_2_2_3_4_1000_in3)
          begin :bnn_N_Mux_2_2_3_4_1000
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1000_out1 = bnn_Minus_2S_2S_4_985_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1000_out1 = bnn_N_Mux_2_2_3_4_1000_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1001
         assign bnn_Add_4Sx3S_4S_1_1001_out1 = bnn_Add_3Sx3S_4S_4_987_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_986_out1[1]}}, bnn_N_Mux_2_2_3_4_986_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_13_mi61 or s_reg_1112 or s_reg_882 or s_reg_997 or bnn_N_Mux_64_2_2_1_1636_out1[34] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1002_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1002_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[34], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1002_in1 = Bline_buffer_13_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1002_in1 = s_reg_997;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1002_in1 = s_reg_882;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1002
         assign bnn_Minus_2S_2S_1_1002_out1 = -bnn_Minus_2S_2S_1_1002_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_12_mi61 or s_reg_1112 or s_reg_877 or s_reg_995 or bnn_N_Mux_64_2_2_1_1636_out1[33] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1003_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1003_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1003_in3 = Bline_buffer_12_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1003_in3 = s_reg_995;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1003_in3 = s_reg_877;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_988_out1 or bnn_N_Mux_2_2_3_1_1003_in3)
          begin :bnn_N_Mux_2_2_3_1_1003
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1003_out1 = bnn_Minus_2S_2S_1_988_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1003_out1 = bnn_N_Mux_2_2_3_1_1003_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1004
         assign bnn_Add_4Sx2S_4S_1_1004_out1 = bnn_Add_3Sx3S_4S_1_990_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_989_out1[1]}}, bnn_N_Mux_2_2_3_1_989_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1005
         assign bnn_Minus_2S_2S_1_1005_out1 = -bnn_Minus_2S_2S_1_1002_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_991_out1 or bnn_N_Mux_2_2_3_1_1003_in3)
          begin :bnn_N_Mux_2_2_3_1_1006
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1006_out1 = bnn_Minus_2S_2S_1_991_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1006_out1 = bnn_N_Mux_2_2_3_1_1003_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1007
         assign bnn_Add_3Sx3S_4S_1_1007_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_993_out1[1]}}, bnn_N_Mux_2_2_3_1_993_out1} + {bnn_Add_2Sx2S_3S_1_992_out1[2], bnn_Add_2Sx2S_3S_1_992_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1008
         assign bnn_Minus_2S_2S_1_1008_out1 = -bnn_Minus_2S_2S_1_1002_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1009
         assign bnn_Add_2Sx2S_3S_1_1009_out1 = {bnn_N_Mux_2_2_3_1_995_out1[1], bnn_N_Mux_2_2_3_1_995_out1} + {bnn_N_Mux_2_2_3_1_994_out1[1], bnn_N_Mux_2_2_3_1_994_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_5_mi61 or s_reg_1112 or s_reg_898 or s_reg_984 or bnn_N_Mux_2_2_3_1_1879_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1010_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1010_in3 = bnn_N_Mux_2_2_3_1_1879_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1010_in3 = Bline_buffer_5_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1010_in3 = s_reg_984;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1010_in3 = s_reg_898;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_996_out1 or bnn_N_Mux_2_2_3_1_1010_in3)
          begin :bnn_N_Mux_2_2_3_1_1010
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1010_out1 = bnn_Minus_2S_2S_1_996_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1010_out1 = bnn_N_Mux_2_2_3_1_1010_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_5_mi61 or s_reg_1112 or s_reg_898 or bnn_N_Mux_2_2_3_1_1879_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1011_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1011_in3 = bnn_N_Mux_2_2_3_1_1879_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1011_in3 = Bline_buffer_5_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1011_in3 = s_reg_898;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_997_out1 or bnn_N_Mux_2_2_3_1_1011_in3)
          begin :bnn_N_Mux_2_2_3_1_1011
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1011_out1 = bnn_Minus_2S_2S_1_997_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1011_out1 = bnn_N_Mux_2_2_3_1_1011_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_4_mi61 or s_reg_1112 or s_reg_888 or bnn_N_Mux_2_2_3_1_1868_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1012_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1012_in3 = bnn_N_Mux_2_2_3_1_1868_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1012_in3 = Bline_buffer_4_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1012_in3 = s_reg_888;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_998_out1 or bnn_N_Mux_2_2_3_1_1012_in3)
          begin :bnn_N_Mux_2_2_3_1_1012
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1012_out1 = bnn_Minus_2S_2S_1_998_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1012_out1 = bnn_N_Mux_2_2_3_1_1012_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_6_mi61 or s_reg_1112 or s_reg_909 or s_reg_998 or bnn_N_Mux_2_2_3_1_1890_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1013_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1013_in1 = bnn_N_Mux_2_2_3_1_1890_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1013_in1 = Bline_buffer_6_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1013_in1 = s_reg_998;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1013_in1 = s_reg_909;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1013
         assign bnn_Minus_2S_2S_1_1013_out1 = -bnn_Minus_2S_2S_1_1013_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_6_mi61 or s_reg_1112 or s_reg_909 or bnn_N_Mux_2_2_3_1_1890_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1014_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1014_in1 = bnn_N_Mux_2_2_3_1_1890_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1014_in1 = Bline_buffer_6_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1014_in1 = s_reg_909;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1014
         assign bnn_Minus_2S_2S_4_1014_out1 = -bnn_Minus_2S_2S_4_1014_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1015
         assign bnn_Minus_2S_2S_4_1015_out1 = -bnn_Minus_2S_2S_1_997_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_999_out1 or bnn_N_Mux_3_2_6_4_957_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1016
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_1016_out1 = bnn_Minus_2S_2S_1_999_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1016_out1 = bnn_N_Mux_3_2_6_4_957_out1_slice;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1017
         assign bnn_Add_4Sx3S_4S_1_1017_out1 = bnn_Add_4Sx3S_4S_1_1001_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1000_out1[1]}}, bnn_N_Mux_2_2_3_4_1000_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_13_mi61 or s_reg_1112 or s_reg_882 or s_reg_997 or bnn_N_Mux_64_2_2_1_1636_out1[34] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1018_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1018_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[34], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1018_in3 = Bline_buffer_13_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1018_in3 = s_reg_997;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1018_in3 = s_reg_882;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1002_out1 or bnn_N_Mux_2_2_3_1_1018_in3)
          begin :bnn_N_Mux_2_2_3_1_1018
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1018_out1 = bnn_Minus_2S_2S_1_1002_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1018_out1 = bnn_N_Mux_2_2_3_1_1018_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1019
         assign bnn_Add_4Sx2S_4S_1_1019_out1 = bnn_Add_4Sx2S_4S_1_1004_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1003_out1[1]}}, bnn_N_Mux_2_2_3_1_1003_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_14_mi61 or s_reg_1112 or s_reg_889 or s_reg_999 or bnn_N_Mux_64_2_2_1_1636_out1[35] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1020_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1020_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1020_in1 = Bline_buffer_14_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1020_in1 = s_reg_999;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1020_in1 = s_reg_889;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1020
         assign bnn_Minus_2S_2S_1_1020_out1 = -bnn_Minus_2S_2S_1_1020_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1005_out1 or bnn_N_Mux_2_2_3_1_1018_in3)
          begin :bnn_N_Mux_2_2_3_1_1021
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1021_out1 = bnn_Minus_2S_2S_1_1005_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1021_out1 = bnn_N_Mux_2_2_3_1_1018_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1022
         assign bnn_Add_4Sx2S_4S_1_1022_out1 = bnn_Add_3Sx3S_4S_1_1007_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1006_out1[1]}}, bnn_N_Mux_2_2_3_1_1006_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1023
         assign bnn_Minus_2S_2S_1_1023_out1 = -bnn_Minus_2S_2S_1_1020_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1008_out1 or bnn_N_Mux_2_2_3_1_1018_in3)
          begin :bnn_N_Mux_2_2_3_1_1024
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1024_out1 = bnn_Minus_2S_2S_1_1008_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1024_out1 = bnn_N_Mux_2_2_3_1_1018_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1025
         assign bnn_Add_3Sx3S_4S_1_1025_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1010_out1[1]}}, bnn_N_Mux_2_2_3_1_1010_out1} + {bnn_Add_2Sx2S_3S_1_1009_out1[2], bnn_Add_2Sx2S_3S_1_1009_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_14_mi61 or s_reg_1112 or s_reg_889 or bnn_N_Mux_64_2_2_1_1636_out1[35] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1026_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1026_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1026_in1 = Bline_buffer_14_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1026_in1 = s_reg_889;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1026
         assign bnn_Minus_2S_2S_4_1026_out1 = -bnn_Minus_2S_2S_4_1026_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1027
         assign bnn_Add_2Sx2S_3S_1_1027_out1 = {bnn_N_Mux_2_2_3_1_1012_out1[1], bnn_N_Mux_2_2_3_1_1012_out1} + {bnn_N_Mux_2_2_3_1_1011_out1[1], bnn_N_Mux_2_2_3_1_1011_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_6_mi61 or s_reg_1112 or s_reg_909 or s_reg_998 or bnn_N_Mux_2_2_3_1_1890_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1028_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1028_in3 = bnn_N_Mux_2_2_3_1_1890_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1028_in3 = Bline_buffer_6_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1028_in3 = s_reg_998;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1028_in3 = s_reg_909;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_976_ctrl1 or bnn_Minus_2S_2S_1_1013_out1 or bnn_N_Mux_2_2_3_1_1028_in3)
          begin :bnn_N_Mux_2_2_3_1_1028
            if (bnn_N_Mux_2_2_3_1_976_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1028_out1 = bnn_Minus_2S_2S_1_1013_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1028_out1 = bnn_N_Mux_2_2_3_1_1028_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_6_mi61 or s_reg_1112 or s_reg_909 or bnn_N_Mux_2_2_3_1_1890_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1029_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1029_in3 = bnn_N_Mux_2_2_3_1_1890_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1029_in3 = Bline_buffer_6_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1029_in3 = s_reg_909;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_Minus_2S_2S_4_1014_out1 or bnn_N_Mux_2_2_3_4_1029_in3)
          begin :bnn_N_Mux_2_2_3_4_1029
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_1029_out1 = bnn_Minus_2S_2S_4_1014_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1029_out1 = bnn_N_Mux_2_2_3_4_1029_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1011_in3 or bnn_Minus_2S_2S_4_1015_out1)
          begin :bnn_N_Mux_2_2_3_4_1030
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1030_out1 = bnn_Minus_2S_2S_4_1015_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1030_out1 = bnn_N_Mux_2_2_3_1_1011_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_7_mi61 or s_reg_1112 or s_reg_917 or s_reg_977 or bnn_N_Mux_2_2_3_1_1901_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1031_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1031_in1 = bnn_N_Mux_2_2_3_1_1901_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1031_in1 = Bline_buffer_7_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1031_in1 = s_reg_977;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1031_in1 = s_reg_917;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1031
         assign bnn_Minus_2S_2S_1_1031_out1 = -bnn_Minus_2S_2S_1_1031_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_7_mi61 or s_reg_1112 or s_reg_917 or bnn_N_Mux_2_2_3_1_1901_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1032_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1032_in1 = bnn_N_Mux_2_2_3_1_1901_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1032_in1 = Bline_buffer_7_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1032_in1 = s_reg_917;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1032
         assign bnn_Minus_2S_2S_1_1032_out1 = -bnn_Minus_2S_2S_1_1032_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1033
         assign bnn_Minus_2S_2S_1_1033_out1 = -bnn_Minus_2S_2S_4_1014_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1034
         assign bnn_Add_4Sx2S_5S_1_1034_out1 = {bnn_Add_4Sx3S_4S_1_1017_out1[3], bnn_Add_4Sx3S_4S_1_1017_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1016_out1[1]}}, bnn_N_Mux_2_2_3_1_1016_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_8_mi61 or s_reg_1112 or s_reg_925 or bnn_N_Mux_2_2_3_1_1912_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1035_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1035_in1 = bnn_N_Mux_2_2_3_1_1912_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1035_in1 = Bline_buffer_8_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1035_in1 = s_reg_925;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1035
         assign bnn_Minus_2S_2S_1_1035_out1 = -bnn_Minus_2S_2S_1_1035_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1036
         assign bnn_Minus_2S_2S_1_1036_out1 = -bnn_Minus_2S_2S_1_1032_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1037
         assign bnn_Add_4Sx2S_5S_1_1037_out1 = {bnn_Add_4Sx2S_4S_1_1019_out1[3], bnn_Add_4Sx2S_4S_1_1019_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1018_out1[1]}}, bnn_N_Mux_2_2_3_1_1018_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_14_mi61 or s_reg_1112 or s_reg_889 or s_reg_999 or bnn_N_Mux_64_2_2_1_1636_out1[35] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1038_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1038_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1038_in3 = Bline_buffer_14_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1038_in3 = s_reg_999;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1038_in3 = s_reg_889;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1020_out1 or bnn_N_Mux_2_2_3_1_1038_in3)
          begin :bnn_N_Mux_2_2_3_1_1038
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1038_out1 = bnn_Minus_2S_2S_1_1020_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1038_out1 = bnn_N_Mux_2_2_3_1_1038_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1039
         assign bnn_Add_4Sx2S_4S_1_1039_out1 = bnn_Add_4Sx2S_4S_1_1022_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1021_out1[1]}}, bnn_N_Mux_2_2_3_1_1021_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_15_mi61 or s_reg_1112 or s_reg_899 or s_reg_996 or bnn_N_Mux_64_2_2_1_1636_out1[36] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1040_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1040_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1040_in1 = Bline_buffer_15_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1040_in1 = s_reg_996;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1040_in1 = s_reg_899;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1040
         assign bnn_Minus_2S_2S_1_1040_out1 = -bnn_Minus_2S_2S_1_1040_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1023_out1 or bnn_N_Mux_2_2_3_1_1038_in3)
          begin :bnn_N_Mux_2_2_3_1_1041
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1041_out1 = bnn_Minus_2S_2S_1_1023_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1041_out1 = bnn_N_Mux_2_2_3_1_1038_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1042
         assign bnn_Add_4Sx2S_4S_1_1042_out1 = bnn_Add_3Sx3S_4S_1_1025_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1024_out1[1]}}, bnn_N_Mux_2_2_3_1_1024_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_15_mi61 or s_reg_1112 or s_reg_899 or bnn_N_Mux_64_2_2_1_1636_out1[36] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1043_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1043_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1043_in1 = Bline_buffer_15_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1043_in1 = s_reg_899;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1043
         assign bnn_Minus_2S_2S_4_1043_out1 = -bnn_Minus_2S_2S_4_1043_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_14_mi61 or s_reg_1112 or s_reg_889 or bnn_N_Mux_64_2_2_1_1636_out1[35] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1044_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1044_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1044_in3 = Bline_buffer_14_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1044_in3 = s_reg_889;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1026_out1 or bnn_N_Mux_2_2_3_4_1044_in3)
          begin :bnn_N_Mux_2_2_3_4_1044
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1044_out1 = bnn_Minus_2S_2S_4_1026_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1044_out1 = bnn_N_Mux_2_2_3_4_1044_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1045
         assign bnn_Add_3Sx3S_4S_4_1045_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1028_out1[1]}}, bnn_N_Mux_2_2_3_1_1028_out1} + {bnn_Add_2Sx2S_3S_1_1027_out1[2], bnn_Add_2Sx2S_3S_1_1027_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1046
         assign bnn_Minus_2S_2S_4_1046_out1 = -bnn_Minus_2S_2S_4_1043_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1047
         assign bnn_Add_2Sx2S_3S_1_1047_out1 = {bnn_N_Mux_2_2_3_4_1030_out1[1], bnn_N_Mux_2_2_3_4_1030_out1} + {bnn_N_Mux_2_2_3_4_1029_out1[1], bnn_N_Mux_2_2_3_4_1029_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_7_mi61 or s_reg_1112 or s_reg_917 or s_reg_977 or bnn_N_Mux_2_2_3_1_1901_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1048_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1048_in3 = bnn_N_Mux_2_2_3_1_1901_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1048_in3 = Bline_buffer_7_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1048_in3 = s_reg_977;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1048_in3 = s_reg_917;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_976_ctrl1 or bnn_Minus_2S_2S_1_1031_out1 or bnn_N_Mux_2_2_3_1_1048_in3)
          begin :bnn_N_Mux_2_2_3_1_1048
            if (bnn_N_Mux_2_2_3_1_976_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1048_out1 = bnn_Minus_2S_2S_1_1031_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1048_out1 = bnn_N_Mux_2_2_3_1_1048_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_7_mi61 or s_reg_1112 or s_reg_917 or bnn_N_Mux_2_2_3_1_1901_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1049_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1049_in3 = bnn_N_Mux_2_2_3_1_1901_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1049_in3 = Bline_buffer_7_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1049_in3 = s_reg_917;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1032_out1 or bnn_N_Mux_2_2_3_1_1049_in3)
          begin :bnn_N_Mux_2_2_3_1_1049
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1049_out1 = bnn_Minus_2S_2S_1_1032_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1049_out1 = bnn_N_Mux_2_2_3_1_1049_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_4_1029_in3 or bnn_Minus_2S_2S_1_1033_out1)
          begin :bnn_N_Mux_2_2_3_1_1050
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1050_out1 = bnn_Minus_2S_2S_1_1033_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1050_out1 = bnn_N_Mux_2_2_3_4_1029_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1051
         assign bnn_Minus_2S_2S_1_1051_out1 = -bnn_Minus_2S_2S_1_1035_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_8_mi61 or s_reg_1112 or s_reg_925 or bnn_N_Mux_2_2_3_1_1912_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1052_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1052_in3 = bnn_N_Mux_2_2_3_1_1912_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1052_in3 = Bline_buffer_8_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1052_in3 = s_reg_925;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1035_out1 or bnn_N_Mux_2_2_3_1_1052_in3)
          begin :bnn_N_Mux_2_2_3_1_1052
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1052_out1 = bnn_Minus_2S_2S_1_1035_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1052_out1 = bnn_N_Mux_2_2_3_1_1052_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1036_out1 or bnn_N_Mux_2_2_3_1_1049_in3)
          begin :bnn_N_Mux_2_2_3_1_1053
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1053_out1 = bnn_Minus_2S_2S_1_1036_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1053_out1 = bnn_N_Mux_2_2_3_1_1049_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_9_mi61 or s_reg_1112 or s_reg_933 or bnn_N_Mux_2_2_3_1_2164_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1054_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1054_in1 = bnn_N_Mux_2_2_3_1_2164_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1054_in1 = Bline_buffer_9_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1054_in1 = s_reg_933;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1054
         assign bnn_Minus_2S_2S_1_1054_out1 = -bnn_Minus_2S_2S_1_1054_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_31_mi61 or s_reg_1112 or s_reg_879 or bnn_N_Mux_2_2_3_1_1933_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1055_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1055_in1 = bnn_N_Mux_2_2_3_1_1933_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1055_in1 = Bline_buffer_31_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1055_in1 = s_reg_879;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1055
         assign bnn_Minus_2S_2S_1_1055_out1 = -bnn_Minus_2S_2S_1_1055_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_30_mi61 or s_reg_1112 or s_reg_891 or bnn_N_Mux_2_2_3_1_2176_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1056_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1056_in1 = bnn_N_Mux_2_2_3_1_2176_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1056_in1 = Bline_buffer_30_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1056_in1 = s_reg_891;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1056
         assign bnn_Minus_2S_2S_1_1056_out1 = -bnn_Minus_2S_2S_1_1056_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1057
         assign bnn_Add_4Sx2S_5S_1_1057_out1 = {bnn_Add_4Sx2S_4S_1_1039_out1[3], bnn_Add_4Sx2S_4S_1_1039_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1038_out1[1]}}, bnn_N_Mux_2_2_3_1_1038_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_15_mi61 or s_reg_1112 or s_reg_899 or s_reg_996 or bnn_N_Mux_64_2_2_1_1636_out1[36] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1058_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1058_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1058_in3 = Bline_buffer_15_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1058_in3 = s_reg_996;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1058_in3 = s_reg_899;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_939 or s_reg_944 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_1058_ctrl1
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_1058_ctrl1 = s_reg_944;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1058_ctrl1 = s_reg_939;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1040_out1 or bnn_N_Mux_2_2_3_1_1058_in3 or bnn_N_Mux_2_2_3_1_1058_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1058
            if (bnn_N_Mux_2_2_3_1_1058_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1058_out1 = bnn_Minus_2S_2S_1_1040_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1058_out1 = bnn_N_Mux_2_2_3_1_1058_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1059
         assign bnn_Add_4Sx2S_4S_1_1059_out1 = bnn_Add_4Sx2S_4S_1_1042_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1041_out1[1]}}, bnn_N_Mux_2_2_3_1_1041_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_16_mi61 or s_reg_1112 or s_reg_910 or bnn_N_Mux_64_2_2_1_1636_out1[37] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1060_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1060_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[37], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1060_in1 = Bline_buffer_16_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1060_in1 = s_reg_910;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1060
         assign bnn_Minus_2S_2S_4_1060_out1 = -bnn_Minus_2S_2S_4_1060_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_15_mi61 or s_reg_1112 or s_reg_899 or bnn_N_Mux_64_2_2_1_1636_out1[36] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1061_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1061_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1061_in3 = Bline_buffer_15_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1061_in3 = s_reg_899;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1043_out1 or bnn_N_Mux_2_2_3_4_1061_in3)
          begin :bnn_N_Mux_2_2_3_4_1061
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1061_out1 = bnn_Minus_2S_2S_4_1043_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1061_out1 = bnn_N_Mux_2_2_3_4_1061_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1062
         assign bnn_Add_4Sx3S_4S_1_1062_out1 = bnn_Add_3Sx3S_4S_4_1045_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1044_out1[1]}}, bnn_N_Mux_2_2_3_4_1044_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1063
         assign bnn_Minus_2S_2S_4_1063_out1 = -bnn_Minus_2S_2S_4_1060_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1046_out1 or bnn_N_Mux_2_2_3_4_1061_in3)
          begin :bnn_N_Mux_2_2_3_4_1064
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1064_out1 = bnn_Minus_2S_2S_4_1046_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1064_out1 = bnn_N_Mux_2_2_3_4_1061_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1065
         assign bnn_Add_3Sx3S_4S_1_1065_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1048_out1[1]}}, bnn_N_Mux_2_2_3_1_1048_out1} + {bnn_Add_2Sx2S_3S_1_1047_out1[2], bnn_Add_2Sx2S_3S_1_1047_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1066
         assign bnn_Minus_2S_2S_4_1066_out1 = -bnn_Minus_2S_2S_4_1060_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1067
         assign bnn_Add_2Sx2S_3S_1_1067_out1 = {bnn_N_Mux_2_2_3_1_1050_out1[1], bnn_N_Mux_2_2_3_1_1050_out1} + {bnn_N_Mux_2_2_3_1_1049_out1[1], bnn_N_Mux_2_2_3_1_1049_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1051_out1 or bnn_N_Mux_2_2_3_1_1052_in3)
          begin :bnn_N_Mux_2_2_3_1_1068
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1068_out1 = bnn_Minus_2S_2S_1_1051_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1068_out1 = bnn_N_Mux_2_2_3_1_1052_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_17_mi61 or s_reg_1112 or s_reg_918 or bnn_N_Mux_64_2_2_1_1636_out1[38] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1069_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1069_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[38], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1069_in1 = Bline_buffer_17_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1069_in1 = s_reg_918;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1069
         assign bnn_Minus_2S_2S_4_1069_out1 = -bnn_Minus_2S_2S_4_1069_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1070
         assign bnn_Add_2Sx2S_3S_1_1070_out1 = {bnn_N_Mux_2_2_3_1_1053_out1[1], bnn_N_Mux_2_2_3_1_1053_out1} + {bnn_N_Mux_2_2_3_1_1052_out1[1], bnn_N_Mux_2_2_3_1_1052_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_9_mi61 or s_reg_1112 or s_reg_933 or bnn_N_Mux_2_2_3_1_2164_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1071_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1071_in3 = bnn_N_Mux_2_2_3_1_2164_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1071_in3 = Bline_buffer_9_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1071_in3 = s_reg_933;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1054_out1 or bnn_N_Mux_2_2_3_1_1071_in3)
          begin :bnn_N_Mux_2_2_3_1_1071
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1071_out1 = bnn_Minus_2S_2S_1_1054_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1071_out1 = bnn_N_Mux_2_2_3_1_1071_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_31_mi61 or s_reg_1112 or s_reg_879 or bnn_N_Mux_2_2_3_1_1933_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1072_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1072_in3 = bnn_N_Mux_2_2_3_1_1933_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1072_in3 = Bline_buffer_31_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1072_in3 = s_reg_879;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1055_out1 or bnn_N_Mux_2_2_3_1_1072_in3)
          begin :bnn_N_Mux_2_2_3_1_1072
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1072_out1 = bnn_Minus_2S_2S_1_1055_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1072_out1 = bnn_N_Mux_2_2_3_1_1072_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_30_mi61 or s_reg_1112 or s_reg_891 or bnn_N_Mux_2_2_3_1_2176_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1073_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1073_in3 = bnn_N_Mux_2_2_3_1_2176_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1073_in3 = Bline_buffer_30_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1073_in3 = s_reg_891;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1056_out1 or bnn_N_Mux_2_2_3_1_1073_in3)
          begin :bnn_N_Mux_2_2_3_1_1073
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1073_out1 = bnn_Minus_2S_2S_1_1056_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1073_out1 = bnn_N_Mux_2_2_3_1_1073_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_32_mi61 or s_reg_1112 or s_reg_880 or bnn_N_Mux_2_2_3_1_1944_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1074_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1074_in1 = bnn_N_Mux_2_2_3_1_1944_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1074_in1 = Bline_buffer_32_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1074_in1 = s_reg_880;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1074
         assign bnn_Minus_2S_2S_1_1074_out1 = -bnn_Minus_2S_2S_1_1074_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1075
         assign bnn_Add_4Sx2S_5S_1_1075_out1 = {bnn_Add_4Sx2S_4S_1_1059_out1[3], bnn_Add_4Sx2S_4S_1_1059_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1058_out1[1]}}, bnn_N_Mux_2_2_3_1_1058_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_16_mi61 or s_reg_1112 or s_reg_910 or bnn_N_Mux_64_2_2_1_1636_out1[37] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1076_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1076_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[37], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1076_in3 = Bline_buffer_16_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1076_in3 = s_reg_910;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1060_out1 or bnn_N_Mux_2_2_3_4_1076_in3)
          begin :bnn_N_Mux_2_2_3_4_1076
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1076_out1 = bnn_Minus_2S_2S_4_1060_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1076_out1 = bnn_N_Mux_2_2_3_4_1076_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1077
         assign bnn_Add_4Sx3S_4S_1_1077_out1 = bnn_Add_4Sx3S_4S_1_1062_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1061_out1[1]}}, bnn_N_Mux_2_2_3_4_1061_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1078
         assign bnn_Minus_2S_2S_4_1078_out1 = -bnn_Minus_2S_2S_4_1069_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1063_out1 or bnn_N_Mux_2_2_3_4_1076_in3)
          begin :bnn_N_Mux_2_2_3_4_1079
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1079_out1 = bnn_Minus_2S_2S_4_1063_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1079_out1 = bnn_N_Mux_2_2_3_4_1076_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1080
         assign bnn_Add_4Sx3S_4S_1_1080_out1 = bnn_Add_3Sx3S_4S_1_1065_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1064_out1[1]}}, bnn_N_Mux_2_2_3_4_1064_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1081
         assign bnn_Minus_2S_2S_4_1081_out1 = -bnn_Minus_2S_2S_4_1069_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1066_out1 or bnn_N_Mux_2_2_3_4_1076_in3)
          begin :bnn_N_Mux_2_2_3_4_1082
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1082_out1 = bnn_Minus_2S_2S_4_1066_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1082_out1 = bnn_N_Mux_2_2_3_4_1076_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1083
         assign bnn_Add_3Sx3S_4S_1_1083_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1068_out1[1]}}, bnn_N_Mux_2_2_3_1_1068_out1} + {bnn_Add_2Sx2S_3S_1_1067_out1[2], bnn_Add_2Sx2S_3S_1_1067_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_32_mi61 or s_reg_1112 or s_reg_880 or s_reg_956 or bnn_N_Mux_2_2_3_1_1944_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1084_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1084_in1 = bnn_N_Mux_2_2_3_1_1944_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1084_in1 = Bline_buffer_32_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1084_in1 = s_reg_956;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1084_in1 = s_reg_880;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1084
         assign bnn_Minus_2S_2S_1_1084_out1 = -bnn_Minus_2S_2S_1_1084_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_31_mi61 or s_reg_1112 or s_reg_879 or s_reg_950 or bnn_N_Mux_2_2_3_1_1933_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1085_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1085_in1 = bnn_N_Mux_2_2_3_1_1933_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1085_in1 = Bline_buffer_31_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1085_in1 = s_reg_950;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1085_in1 = s_reg_879;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1085
         assign bnn_Minus_2S_2S_1_1085_out1 = -bnn_Minus_2S_2S_1_1085_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_18_mi61 or s_reg_1112 or s_reg_926 or bnn_N_Mux_64_2_2_1_1636_out1[39] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1086_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1086_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[39], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1086_in1 = Bline_buffer_18_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1086_in1 = s_reg_926;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1086
         assign bnn_Minus_2S_2S_4_1086_out1 = -bnn_Minus_2S_2S_4_1086_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_17_mi61 or s_reg_1112 or s_reg_918 or bnn_N_Mux_64_2_2_1_1636_out1[38] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1087_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1087_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[38], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1087_in3 = Bline_buffer_17_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1087_in3 = s_reg_918;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1069_out1 or bnn_N_Mux_2_2_3_4_1087_in3)
          begin :bnn_N_Mux_2_2_3_4_1087
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1087_out1 = bnn_Minus_2S_2S_4_1069_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1087_out1 = bnn_N_Mux_2_2_3_4_1087_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1088
         assign bnn_Add_3Sx3S_4S_1_1088_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1071_out1[1]}}, bnn_N_Mux_2_2_3_1_1071_out1} + {bnn_Add_2Sx2S_3S_1_1070_out1[2], bnn_Add_2Sx2S_3S_1_1070_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_40_mi61 or s_reg_1112 or s_reg_902 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1638_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_1089_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1089_in1 = bnn_N_Mux_3_2_6_4_1638_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_1089_in1 = Bline_buffer_40_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1089_in1 = s_reg_902;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1089
         assign bnn_Minus_2S_2S_4_1089_out1 = -bnn_Minus_2S_2S_4_1089_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1090
         assign bnn_Add_2Sx2S_3S_1_1090_out1 = {bnn_N_Mux_2_2_3_1_1073_out1[1], bnn_N_Mux_2_2_3_1_1073_out1} + {bnn_N_Mux_2_2_3_1_1072_out1[1], bnn_N_Mux_2_2_3_1_1072_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_32_mi61 or s_reg_1112 or s_reg_880 or bnn_N_Mux_2_2_3_1_1944_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1091_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1091_in3 = bnn_N_Mux_2_2_3_1_1944_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1091_in3 = Bline_buffer_32_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1091_in3 = s_reg_880;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1074_out1 or bnn_N_Mux_2_2_3_1_1091_in3)
          begin :bnn_N_Mux_2_2_3_1_1091
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1091_out1 = bnn_Minus_2S_2S_1_1074_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1091_out1 = bnn_N_Mux_2_2_3_1_1091_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1092
         assign bnn_Add_4Sx2S_5S_1_1092_out1 = {bnn_Add_4Sx3S_4S_1_1077_out1[3], bnn_Add_4Sx3S_4S_1_1077_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1076_out1[1]}}, bnn_N_Mux_2_2_3_4_1076_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1078_out1 or bnn_N_Mux_2_2_3_4_1087_in3)
          begin :bnn_N_Mux_2_2_3_4_1093
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1093_out1 = bnn_Minus_2S_2S_4_1078_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1093_out1 = bnn_N_Mux_2_2_3_4_1087_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1094
         assign bnn_Add_4Sx3S_4S_1_1094_out1 = bnn_Add_4Sx3S_4S_1_1080_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1079_out1[1]}}, bnn_N_Mux_2_2_3_4_1079_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1095
         assign bnn_Minus_2S_2S_4_1095_out1 = -bnn_Minus_2S_2S_4_1086_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1081_out1 or bnn_N_Mux_2_2_3_4_1087_in3)
          begin :bnn_N_Mux_2_2_3_4_1096
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1096_out1 = bnn_Minus_2S_2S_4_1081_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1096_out1 = bnn_N_Mux_2_2_3_4_1087_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1097
         assign bnn_Add_4Sx2S_4S_1_1097_out1 = bnn_Add_3Sx3S_4S_1_1083_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1082_out1[1]}}, bnn_N_Mux_2_2_3_4_1082_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_32_mi61 or s_reg_1112 or s_reg_880 or s_reg_956 or bnn_N_Mux_2_2_3_1_1944_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1098_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1098_in3 = bnn_N_Mux_2_2_3_1_1944_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1098_in3 = Bline_buffer_32_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1098_in3 = s_reg_956;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1098_in3 = s_reg_880;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1084_out1 or bnn_N_Mux_2_2_3_1_1098_in3)
          begin :bnn_N_Mux_2_2_3_1_1098
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1098_out1 = bnn_Minus_2S_2S_1_1084_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1098_out1 = bnn_N_Mux_2_2_3_1_1098_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_31_mi61 or s_reg_1112 or s_reg_879 or s_reg_950 or bnn_N_Mux_2_2_3_1_1933_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1099_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1099_in3 = bnn_N_Mux_2_2_3_1_1933_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1099_in3 = Bline_buffer_31_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1099_in3 = s_reg_950;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1099_in3 = s_reg_879;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1085_out1 or bnn_N_Mux_2_2_3_1_1099_in3)
          begin :bnn_N_Mux_2_2_3_1_1099
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1099_out1 = bnn_Minus_2S_2S_1_1085_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1099_out1 = bnn_N_Mux_2_2_3_1_1099_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_33_mi61 or s_reg_1112 or s_reg_885 or s_reg_960 or bnn_N_Mux_2_2_3_1_1955_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1100_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1100_in1 = bnn_N_Mux_2_2_3_1_1955_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1100_in1 = Bline_buffer_33_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1100_in1 = s_reg_960;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1100_in1 = s_reg_885;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1100
         assign bnn_Minus_2S_2S_1_1100_out1 = -bnn_Minus_2S_2S_1_1100_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1101
         assign bnn_Minus_2S_2S_1_1101_out1 = -bnn_Minus_2S_2S_1_1100_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1102
         assign bnn_Minus_2S_2S_1_1102_out1 = -bnn_Minus_2S_2S_1_1084_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_19_mi61 or s_reg_1112 or s_reg_934 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1637_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_1103_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1103_in1 = bnn_N_Mux_3_2_6_4_1637_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_1103_in1 = Bline_buffer_19_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1103_in1 = s_reg_934;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1103
         assign bnn_Minus_2S_2S_4_1103_out1 = -bnn_Minus_2S_2S_4_1103_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_18_mi61 or s_reg_1112 or s_reg_926 or bnn_N_Mux_64_2_2_1_1636_out1[39] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1104_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1104_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[39], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1104_in3 = Bline_buffer_18_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1104_in3 = s_reg_926;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1086_out1 or bnn_N_Mux_2_2_3_4_1104_in3)
          begin :bnn_N_Mux_2_2_3_4_1104
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1104_out1 = bnn_Minus_2S_2S_4_1086_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1104_out1 = bnn_N_Mux_2_2_3_4_1104_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1105
         assign bnn_Add_4Sx2S_4S_1_1105_out1 = bnn_Add_3Sx3S_4S_1_1088_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1087_out1[1]}}, bnn_N_Mux_2_2_3_4_1087_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_41_mi61 or s_reg_1112 or s_reg_893 or bnn_N_Mux_64_2_2_1_1636_out1[40] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1106_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1106_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1106_in1 = Bline_buffer_41_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1106_in1 = s_reg_893;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1106
         assign bnn_Minus_2S_2S_4_1106_out1 = -bnn_Minus_2S_2S_4_1106_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_40_mi61 or s_reg_1112 or s_reg_902 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1638_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_1107_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1107_in3 = bnn_N_Mux_3_2_6_4_1638_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1107_in3 = Bline_buffer_40_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1107_in3 = s_reg_902;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1089_out1 or bnn_N_Mux_2_2_3_4_1107_in3)
          begin :bnn_N_Mux_2_2_3_4_1107
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1107_out1 = bnn_Minus_2S_2S_4_1089_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1107_out1 = bnn_N_Mux_2_2_3_4_1107_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1108
         assign bnn_Add_3Sx3S_4S_1_1108_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1091_out1[1]}}, bnn_N_Mux_2_2_3_1_1091_out1} + {bnn_Add_2Sx2S_3S_1_1090_out1[2], bnn_Add_2Sx2S_3S_1_1090_out1};

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1109
         assign bnn_Add_4Sx2S_5S_4_1109_out1 = {bnn_Add_4Sx3S_4S_1_1094_out1[3], bnn_Add_4Sx3S_4S_1_1094_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1093_out1[1]}}, bnn_N_Mux_2_2_3_4_1093_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1095_out1 or bnn_N_Mux_2_2_3_4_1104_in3)
          begin :bnn_N_Mux_2_2_3_4_1110
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1110_out1 = bnn_Minus_2S_2S_4_1095_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1110_out1 = bnn_N_Mux_2_2_3_4_1104_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1111
         assign bnn_Add_4Sx2S_4S_1_1111_out1 = bnn_Add_4Sx2S_4S_1_1097_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1096_out1[1]}}, bnn_N_Mux_2_2_3_4_1096_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_41_mi61 or s_reg_1112 or s_reg_893 or s_reg_981 or bnn_N_Mux_64_2_2_1_1636_out1[40] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1112_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1112_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1112_in1 = Bline_buffer_41_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1112_in1 = s_reg_981;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1112_in1 = s_reg_893;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1112
         assign bnn_Minus_2S_2S_1_1112_out1 = -bnn_Minus_2S_2S_1_1112_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1113
         assign bnn_Add_2Sx2S_3S_1_1113_out1 = {bnn_N_Mux_2_2_3_1_1099_out1[1], bnn_N_Mux_2_2_3_1_1099_out1} + {bnn_N_Mux_2_2_3_1_1098_out1[1], bnn_N_Mux_2_2_3_1_1098_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_33_mi61 or s_reg_1112 or s_reg_885 or s_reg_960 or bnn_N_Mux_2_2_3_1_1955_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1114_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1114_in3 = bnn_N_Mux_2_2_3_1_1955_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1114_in3 = Bline_buffer_33_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1114_in3 = s_reg_960;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1114_in3 = s_reg_885;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1100_out1 or bnn_N_Mux_2_2_3_1_1114_in3)
          begin :bnn_N_Mux_2_2_3_1_1114
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1114_out1 = bnn_Minus_2S_2S_1_1100_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1114_out1 = bnn_N_Mux_2_2_3_1_1114_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1101_out1 or bnn_N_Mux_2_2_3_1_1114_in3)
          begin :bnn_N_Mux_2_2_3_1_1115
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1115_out1 = bnn_Minus_2S_2S_1_1101_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1115_out1 = bnn_N_Mux_2_2_3_1_1114_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1098_in3 or bnn_Minus_2S_2S_1_1102_out1)
          begin :bnn_N_Mux_2_2_3_1_1116
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1116_out1 = bnn_Minus_2S_2S_1_1102_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1116_out1 = bnn_N_Mux_2_2_3_1_1098_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_34_mi61 or s_reg_1112 or s_reg_892 or s_reg_963 or bnn_N_Mux_2_2_3_1_1966_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1117_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1117_in1 = bnn_N_Mux_2_2_3_1_1966_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1117_in1 = Bline_buffer_34_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1117_in1 = s_reg_963;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1117_in1 = s_reg_892;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1117
         assign bnn_Minus_2S_2S_1_1117_out1 = -bnn_Minus_2S_2S_1_1117_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1118
         assign bnn_Minus_2S_2S_1_1118_out1 = -bnn_Minus_2S_2S_1_1117_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1119
         assign bnn_Minus_2S_2S_1_1119_out1 = -bnn_Minus_2S_2S_1_1100_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_19_mi61 or s_reg_1112 or s_reg_934 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1637_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_1120_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1120_in3 = bnn_N_Mux_3_2_6_4_1637_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1120_in3 = Bline_buffer_19_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1120_in3 = s_reg_934;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1103_out1 or bnn_N_Mux_2_2_3_4_1120_in3)
          begin :bnn_N_Mux_2_2_3_4_1120
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1120_out1 = bnn_Minus_2S_2S_4_1103_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1120_out1 = bnn_N_Mux_2_2_3_4_1120_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1121
         assign bnn_Add_4Sx2S_4S_1_1121_out1 = bnn_Add_4Sx2S_4S_1_1105_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1104_out1[1]}}, bnn_N_Mux_2_2_3_4_1104_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_42_mi61 or s_reg_1112 or s_reg_903 or bnn_N_Mux_64_2_2_1_1636_out1[41] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1122_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1122_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1122_in1 = Bline_buffer_42_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1122_in1 = s_reg_903;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1122
         assign bnn_Minus_2S_2S_4_1122_out1 = -bnn_Minus_2S_2S_4_1122_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_41_mi61 or s_reg_1112 or s_reg_893 or bnn_N_Mux_64_2_2_1_1636_out1[40] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1123_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1123_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1123_in3 = Bline_buffer_41_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1123_in3 = s_reg_893;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1106_out1 or bnn_N_Mux_2_2_3_4_1123_in3)
          begin :bnn_N_Mux_2_2_3_4_1123
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1123_out1 = bnn_Minus_2S_2S_4_1106_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1123_out1 = bnn_N_Mux_2_2_3_4_1123_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1124
         assign bnn_Add_4Sx2S_4S_1_1124_out1 = bnn_Add_3Sx3S_4S_1_1108_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1107_out1[1]}}, bnn_N_Mux_2_2_3_4_1107_out1};

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1125
         assign bnn_Add_4Sx2S_5S_1_1125_out1 = {bnn_Add_4Sx2S_4S_1_1111_out1[3], bnn_Add_4Sx2S_4S_1_1111_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1110_out1[1]}}, bnn_N_Mux_2_2_3_4_1110_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_42_mi61 or s_reg_1112 or s_reg_903 or s_reg_985 or bnn_N_Mux_64_2_2_1_1636_out1[41] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1126_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1126_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1126_in1 = Bline_buffer_42_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1126_in1 = s_reg_985;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1126_in1 = s_reg_903;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1126
         assign bnn_Minus_2S_2S_1_1126_out1 = -bnn_Minus_2S_2S_1_1126_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_41_mi61 or s_reg_1112 or s_reg_893 or s_reg_981 or bnn_N_Mux_64_2_2_1_1636_out1[40] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1127_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1127_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1127_in3 = Bline_buffer_41_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1127_in3 = s_reg_981;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1127_in3 = s_reg_893;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1112_out1 or bnn_N_Mux_2_2_3_1_1127_in3)
          begin :bnn_N_Mux_2_2_3_1_1127
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1127_out1 = bnn_Minus_2S_2S_1_1112_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1127_out1 = bnn_N_Mux_2_2_3_1_1127_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1128
         assign bnn_Add_3Sx3S_4S_1_1128_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1114_out1[1]}}, bnn_N_Mux_2_2_3_1_1114_out1} + {bnn_Add_2Sx2S_3S_1_1113_out1[2], bnn_Add_2Sx2S_3S_1_1113_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1129
         assign bnn_Minus_2S_2S_1_1129_out1 = -bnn_Minus_2S_2S_1_1126_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1130
         assign bnn_Add_2Sx2S_3S_1_1130_out1 = {bnn_N_Mux_2_2_3_1_1116_out1[1], bnn_N_Mux_2_2_3_1_1116_out1} + {bnn_N_Mux_2_2_3_1_1115_out1[1], bnn_N_Mux_2_2_3_1_1115_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_34_mi61 or s_reg_1112 or s_reg_892 or s_reg_963 or bnn_N_Mux_2_2_3_1_1966_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1131_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1131_in3 = bnn_N_Mux_2_2_3_1_1966_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1131_in3 = Bline_buffer_34_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1131_in3 = s_reg_963;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1131_in3 = s_reg_892;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1117_out1 or bnn_N_Mux_2_2_3_1_1131_in3)
          begin :bnn_N_Mux_2_2_3_1_1131
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1131_out1 = bnn_Minus_2S_2S_1_1117_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1131_out1 = bnn_N_Mux_2_2_3_1_1131_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1118_out1 or bnn_N_Mux_2_2_3_1_1131_in3)
          begin :bnn_N_Mux_2_2_3_1_1132
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1132_out1 = bnn_Minus_2S_2S_1_1118_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1132_out1 = bnn_N_Mux_2_2_3_1_1131_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1114_in3 or bnn_Minus_2S_2S_1_1119_out1)
          begin :bnn_N_Mux_2_2_3_1_1133
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1133_out1 = bnn_Minus_2S_2S_1_1119_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1133_out1 = bnn_N_Mux_2_2_3_1_1114_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_35_mi61 or s_reg_1112 or s_reg_901 or s_reg_966 or bnn_N_Mux_2_2_3_1_1977_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1134_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1134_in1 = bnn_N_Mux_2_2_3_1_1977_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1134_in1 = Bline_buffer_35_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1134_in1 = s_reg_966;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1134_in1 = s_reg_901;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1134
         assign bnn_Minus_2S_2S_1_1134_out1 = -bnn_Minus_2S_2S_1_1134_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1135
         assign bnn_Minus_2S_2S_1_1135_out1 = -bnn_Minus_2S_2S_1_1134_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1136
         assign bnn_Minus_2S_2S_1_1136_out1 = -bnn_Minus_2S_2S_1_1117_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1137
         assign bnn_Add_4Sx2S_5S_1_1137_out1 = {bnn_Add_4Sx2S_4S_1_1121_out1[3], bnn_Add_4Sx2S_4S_1_1121_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1120_out1[1]}}, bnn_N_Mux_2_2_3_4_1120_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_42_mi61 or s_reg_1112 or s_reg_903 or bnn_N_Mux_64_2_2_1_1636_out1[41] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1138_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1138_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1138_in3 = Bline_buffer_42_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1138_in3 = s_reg_903;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1122_out1 or bnn_N_Mux_2_2_3_4_1138_in3)
          begin :bnn_N_Mux_2_2_3_4_1138
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1138_out1 = bnn_Minus_2S_2S_4_1122_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1138_out1 = bnn_N_Mux_2_2_3_4_1138_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1139
         assign bnn_Add_4Sx2S_4S_1_1139_out1 = bnn_Add_4Sx2S_4S_1_1124_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1123_out1[1]}}, bnn_N_Mux_2_2_3_4_1123_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_43_mi61 or s_reg_1112 or s_reg_913 or s_reg_987 or bnn_N_Mux_64_2_2_1_1636_out1[42] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_4_1140_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_4_1140_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[42], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_4_1140_in1 = Bline_buffer_43_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_4_1140_in1 = s_reg_987;
               end
               
               default: begin
                  bnn_Minus_2S_2S_4_1140_in1 = s_reg_913;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1140
         assign bnn_Minus_2S_2S_4_1140_out1 = -bnn_Minus_2S_2S_4_1140_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_42_mi61 or s_reg_1112 or s_reg_903 or s_reg_985 or bnn_N_Mux_64_2_2_1_1636_out1[41] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1141_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1141_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1141_in3 = Bline_buffer_42_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1141_in3 = s_reg_985;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1141_in3 = s_reg_903;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1126_out1 or bnn_N_Mux_2_2_3_1_1141_in3)
          begin :bnn_N_Mux_2_2_3_1_1141
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1141_out1 = bnn_Minus_2S_2S_1_1126_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1141_out1 = bnn_N_Mux_2_2_3_1_1141_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1142
         assign bnn_Add_4Sx2S_4S_1_1142_out1 = bnn_Add_3Sx3S_4S_1_1128_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1127_out1[1]}}, bnn_N_Mux_2_2_3_1_1127_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1143
         assign bnn_Minus_2S_2S_1_1143_out1 = -bnn_Minus_2S_2S_4_1140_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1129_out1 or bnn_N_Mux_2_2_3_1_1141_in3)
          begin :bnn_N_Mux_2_2_3_1_1144
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1144_out1 = bnn_Minus_2S_2S_1_1129_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1144_out1 = bnn_N_Mux_2_2_3_1_1141_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1145
         assign bnn_Add_3Sx3S_4S_1_1145_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1131_out1[1]}}, bnn_N_Mux_2_2_3_1_1131_out1} + {bnn_Add_2Sx2S_3S_1_1130_out1[2], bnn_Add_2Sx2S_3S_1_1130_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1146
         assign bnn_Minus_2S_2S_1_1146_out1 = -bnn_Minus_2S_2S_4_1140_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1147
         assign bnn_Add_2Sx2S_3S_1_1147_out1 = {bnn_N_Mux_2_2_3_1_1133_out1[1], bnn_N_Mux_2_2_3_1_1133_out1} + {bnn_N_Mux_2_2_3_1_1132_out1[1], bnn_N_Mux_2_2_3_1_1132_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_35_mi61 or s_reg_1112 or s_reg_901 or s_reg_966 or bnn_N_Mux_2_2_3_1_1977_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1148_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1148_in3 = bnn_N_Mux_2_2_3_1_1977_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1148_in3 = Bline_buffer_35_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1148_in3 = s_reg_966;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1148_in3 = s_reg_901;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1134_out1 or bnn_N_Mux_2_2_3_1_1148_in3)
          begin :bnn_N_Mux_2_2_3_1_1148
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1148_out1 = bnn_Minus_2S_2S_1_1134_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1148_out1 = bnn_N_Mux_2_2_3_1_1148_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1135_out1 or bnn_N_Mux_2_2_3_1_1148_in3)
          begin :bnn_N_Mux_2_2_3_1_1149
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1149_out1 = bnn_Minus_2S_2S_1_1135_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1149_out1 = bnn_N_Mux_2_2_3_1_1148_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1131_in3 or bnn_Minus_2S_2S_1_1136_out1)
          begin :bnn_N_Mux_2_2_3_1_1150
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1150_out1 = bnn_Minus_2S_2S_1_1136_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1150_out1 = bnn_N_Mux_2_2_3_1_1131_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_36_mi61 or s_reg_1112 or s_reg_912 or s_reg_969 or bnn_N_Mux_2_2_3_1_1988_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1151_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1151_in1 = bnn_N_Mux_2_2_3_1_1988_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1151_in1 = Bline_buffer_36_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1151_in1 = s_reg_969;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1151_in1 = s_reg_912;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1151
         assign bnn_Minus_2S_2S_1_1151_out1 = -bnn_Minus_2S_2S_1_1151_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1152
         assign bnn_Minus_2S_2S_1_1152_out1 = -bnn_Minus_2S_2S_1_1151_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1153
         assign bnn_Minus_2S_2S_1_1153_out1 = -bnn_Minus_2S_2S_1_1134_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1154
         assign bnn_Add_4Sx2S_5S_1_1154_out1 = {bnn_Add_4Sx2S_4S_1_1139_out1[3], bnn_Add_4Sx2S_4S_1_1139_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1138_out1[1]}}, bnn_N_Mux_2_2_3_4_1138_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_43_mi61 or s_reg_1112 or s_reg_913 or s_reg_987 or bnn_N_Mux_64_2_2_1_1636_out1[42] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_4_1155_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_4_1155_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[42], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_4_1155_in3 = Bline_buffer_43_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_4_1155_in3 = s_reg_987;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_4_1155_in3 = s_reg_913;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1140_out1 or bnn_N_Mux_2_2_3_4_1155_in3)
          begin :bnn_N_Mux_2_2_3_4_1155
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1155_out1 = bnn_Minus_2S_2S_4_1140_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1155_out1 = bnn_N_Mux_2_2_3_4_1155_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1156
         assign bnn_Add_4Sx2S_4S_1_1156_out1 = bnn_Add_4Sx2S_4S_1_1142_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1141_out1[1]}}, bnn_N_Mux_2_2_3_1_1141_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_44_mi61 or s_reg_1112 or s_reg_921 or s_reg_989 or bnn_N_Mux_64_2_2_1_1636_out1[43] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1157_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1157_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[43], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1157_in1 = Bline_buffer_44_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1157_in1 = s_reg_989;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1157_in1 = s_reg_921;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1157
         assign bnn_Minus_2S_2S_1_1157_out1 = -bnn_Minus_2S_2S_1_1157_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1143_out1 or bnn_N_Mux_2_2_3_4_1155_in3)
          begin :bnn_N_Mux_2_2_3_1_1158
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1158_out1 = bnn_Minus_2S_2S_1_1143_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1158_out1 = bnn_N_Mux_2_2_3_4_1155_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1159
         assign bnn_Add_4Sx2S_4S_1_1159_out1 = bnn_Add_3Sx3S_4S_1_1145_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1144_out1[1]}}, bnn_N_Mux_2_2_3_1_1144_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1160
         assign bnn_Minus_2S_2S_1_1160_out1 = -bnn_Minus_2S_2S_1_1157_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1146_out1 or bnn_N_Mux_2_2_3_4_1155_in3)
          begin :bnn_N_Mux_2_2_3_1_1161
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1161_out1 = bnn_Minus_2S_2S_1_1146_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1161_out1 = bnn_N_Mux_2_2_3_4_1155_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1162
         assign bnn_Add_3Sx3S_4S_1_1162_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1148_out1[1]}}, bnn_N_Mux_2_2_3_1_1148_out1} + {bnn_Add_2Sx2S_3S_1_1147_out1[2], bnn_Add_2Sx2S_3S_1_1147_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1163
         assign bnn_Minus_2S_2S_1_1163_out1 = -bnn_Minus_2S_2S_1_1157_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1164
         assign bnn_Add_2Sx2S_3S_1_1164_out1 = {bnn_N_Mux_2_2_3_1_1150_out1[1], bnn_N_Mux_2_2_3_1_1150_out1} + {bnn_N_Mux_2_2_3_1_1149_out1[1], bnn_N_Mux_2_2_3_1_1149_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_36_mi61 or s_reg_1112 or s_reg_912 or s_reg_969 or bnn_N_Mux_2_2_3_1_1988_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1165_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1165_in3 = bnn_N_Mux_2_2_3_1_1988_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1165_in3 = Bline_buffer_36_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1165_in3 = s_reg_969;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1165_in3 = s_reg_912;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1151_out1 or bnn_N_Mux_2_2_3_1_1165_in3)
          begin :bnn_N_Mux_2_2_3_1_1165
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1165_out1 = bnn_Minus_2S_2S_1_1151_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1165_out1 = bnn_N_Mux_2_2_3_1_1165_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1152_out1 or bnn_N_Mux_2_2_3_1_1165_in3)
          begin :bnn_N_Mux_2_2_3_1_1166
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1166_out1 = bnn_Minus_2S_2S_1_1152_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1166_out1 = bnn_N_Mux_2_2_3_1_1165_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1148_in3 or bnn_Minus_2S_2S_1_1153_out1)
          begin :bnn_N_Mux_2_2_3_1_1167
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1167_out1 = bnn_Minus_2S_2S_1_1153_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1167_out1 = bnn_N_Mux_2_2_3_1_1148_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_37_mi61 or s_reg_1112 or s_reg_920 or s_reg_972 or bnn_N_Mux_2_2_3_1_1999_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1168_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1168_in1 = bnn_N_Mux_2_2_3_1_1999_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1168_in1 = Bline_buffer_37_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1168_in1 = s_reg_972;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1168_in1 = s_reg_920;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1168
         assign bnn_Minus_2S_2S_1_1168_out1 = -bnn_Minus_2S_2S_1_1168_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_37_mi61 or s_reg_1112 or s_reg_920 or bnn_N_Mux_2_2_3_1_1999_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1169_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1169_in1 = bnn_N_Mux_2_2_3_1_1999_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1169_in1 = Bline_buffer_37_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1169_in1 = s_reg_920;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1169
         assign bnn_Minus_2S_2S_1_1169_out1 = -bnn_Minus_2S_2S_1_1169_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_36_mi61 or s_reg_1112 or s_reg_912 or bnn_N_Mux_2_2_3_1_1988_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1170_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1170_in1 = bnn_N_Mux_2_2_3_1_1988_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1170_in1 = Bline_buffer_36_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1170_in1 = s_reg_912;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1170
         assign bnn_Minus_2S_2S_1_1170_out1 = -bnn_Minus_2S_2S_1_1170_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_38_mi61 or s_reg_1112 or s_reg_928 or bnn_N_Mux_2_2_3_1_2010_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1171_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1171_in1 = bnn_N_Mux_2_2_3_1_2010_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1171_in1 = Bline_buffer_38_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1171_in1 = s_reg_928;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1171
         assign bnn_Minus_2S_2S_1_1171_out1 = -bnn_Minus_2S_2S_1_1171_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1172
         assign bnn_Minus_2S_2S_1_1172_out1 = -bnn_Minus_2S_2S_1_1169_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1173
         assign bnn_Add_4Sx2S_5S_1_1173_out1 = {bnn_Add_4Sx2S_4S_1_1156_out1[3], bnn_Add_4Sx2S_4S_1_1156_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1155_out1[1]}}, bnn_N_Mux_2_2_3_4_1155_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_44_mi61 or s_reg_1112 or s_reg_921 or s_reg_989 or bnn_N_Mux_64_2_2_1_1636_out1[43] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1174_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1174_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[43], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1174_in3 = Bline_buffer_44_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1174_in3 = s_reg_989;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1174_in3 = s_reg_921;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1157_out1 or bnn_N_Mux_2_2_3_1_1174_in3)
          begin :bnn_N_Mux_2_2_3_1_1174
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1174_out1 = bnn_Minus_2S_2S_1_1157_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1174_out1 = bnn_N_Mux_2_2_3_1_1174_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1175
         assign bnn_Add_4Sx2S_4S_1_1175_out1 = bnn_Add_4Sx2S_4S_1_1159_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1158_out1[1]}}, bnn_N_Mux_2_2_3_1_1158_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_45_mi61 or s_reg_1112 or s_reg_929 or s_reg_991 or bnn_N_Mux_64_2_2_1_1636_out1[44] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1176_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1176_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[44], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1176_in1 = Bline_buffer_45_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1176_in1 = s_reg_991;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1176_in1 = s_reg_929;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1176
         assign bnn_Minus_2S_2S_1_1176_out1 = -bnn_Minus_2S_2S_1_1176_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1160_out1 or bnn_N_Mux_2_2_3_1_1174_in3)
          begin :bnn_N_Mux_2_2_3_1_1177
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1177_out1 = bnn_Minus_2S_2S_1_1160_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1177_out1 = bnn_N_Mux_2_2_3_1_1174_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1178
         assign bnn_Add_4Sx2S_4S_1_1178_out1 = bnn_Add_3Sx3S_4S_1_1162_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1161_out1[1]}}, bnn_N_Mux_2_2_3_1_1161_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1179
         assign bnn_Minus_2S_2S_1_1179_out1 = -bnn_Minus_2S_2S_1_1176_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1163_out1 or bnn_N_Mux_2_2_3_1_1174_in3)
          begin :bnn_N_Mux_2_2_3_1_1180
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1180_out1 = bnn_Minus_2S_2S_1_1163_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1180_out1 = bnn_N_Mux_2_2_3_1_1174_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1181
         assign bnn_Add_3Sx3S_4S_1_1181_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1165_out1[1]}}, bnn_N_Mux_2_2_3_1_1165_out1} + {bnn_Add_2Sx2S_3S_1_1164_out1[2], bnn_Add_2Sx2S_3S_1_1164_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1182
         assign bnn_Minus_2S_2S_1_1182_out1 = -bnn_Minus_2S_2S_1_1176_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1183
         assign bnn_Add_2Sx2S_3S_1_1183_out1 = {bnn_N_Mux_2_2_3_1_1167_out1[1], bnn_N_Mux_2_2_3_1_1167_out1} + {bnn_N_Mux_2_2_3_1_1166_out1[1], bnn_N_Mux_2_2_3_1_1166_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_37_mi61 or s_reg_1112 or s_reg_920 or s_reg_972 or bnn_N_Mux_2_2_3_1_1999_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1184_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1184_in3 = bnn_N_Mux_2_2_3_1_1999_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1184_in3 = Bline_buffer_37_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1184_in3 = s_reg_972;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1184_in3 = s_reg_920;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1168_out1 or bnn_N_Mux_2_2_3_1_1184_in3)
          begin :bnn_N_Mux_2_2_3_1_1184
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1184_out1 = bnn_Minus_2S_2S_1_1168_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1184_out1 = bnn_N_Mux_2_2_3_1_1184_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_37_mi61 or s_reg_1112 or s_reg_920 or bnn_N_Mux_2_2_3_1_1999_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1185_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1185_in3 = bnn_N_Mux_2_2_3_1_1999_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1185_in3 = Bline_buffer_37_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1185_in3 = s_reg_920;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1169_out1 or bnn_N_Mux_2_2_3_1_1185_in3)
          begin :bnn_N_Mux_2_2_3_1_1185
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1185_out1 = bnn_Minus_2S_2S_1_1169_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1185_out1 = bnn_N_Mux_2_2_3_1_1185_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_36_mi61 or s_reg_1112 or s_reg_912 or bnn_N_Mux_2_2_3_1_1988_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1186_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1186_in3 = bnn_N_Mux_2_2_3_1_1988_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1186_in3 = Bline_buffer_36_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1186_in3 = s_reg_912;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1170_out1 or bnn_N_Mux_2_2_3_1_1186_in3)
          begin :bnn_N_Mux_2_2_3_1_1186
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1186_out1 = bnn_Minus_2S_2S_1_1170_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1186_out1 = bnn_N_Mux_2_2_3_1_1186_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1187
         assign bnn_Minus_2S_2S_1_1187_out1 = -bnn_Minus_2S_2S_1_1171_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_38_mi61 or s_reg_1112 or s_reg_928 or bnn_N_Mux_2_2_3_1_2010_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1188_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1188_in3 = bnn_N_Mux_2_2_3_1_2010_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1188_in3 = Bline_buffer_38_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1188_in3 = s_reg_928;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1171_out1 or bnn_N_Mux_2_2_3_1_1188_in3)
          begin :bnn_N_Mux_2_2_3_1_1188
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1188_out1 = bnn_Minus_2S_2S_1_1171_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1188_out1 = bnn_N_Mux_2_2_3_1_1188_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1172_out1 or bnn_N_Mux_2_2_3_1_1185_in3)
          begin :bnn_N_Mux_2_2_3_1_1189
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1189_out1 = bnn_Minus_2S_2S_1_1172_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1189_out1 = bnn_N_Mux_2_2_3_1_1185_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_39_mi61 or s_reg_1112 or s_reg_935 or bnn_N_Mux_2_2_3_1_2190_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1190_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1190_in1 = bnn_N_Mux_2_2_3_1_2190_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1190_in1 = Bline_buffer_39_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1190_in1 = s_reg_935;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1190
         assign bnn_Minus_2S_2S_1_1190_out1 = -bnn_Minus_2S_2S_1_1190_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_61_mi61 or s_reg_1112 or s_reg_896 or bnn_N_Mux_2_2_3_1_2021_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1191_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1191_in1 = bnn_N_Mux_2_2_3_1_2021_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1191_in1 = Bline_buffer_61_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1191_in1 = s_reg_896;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1191
         assign bnn_Minus_2S_2S_1_1191_out1 = -bnn_Minus_2S_2S_1_1191_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_60_mi61 or s_reg_1112 or s_reg_905 or bnn_N_Mux_2_2_3_1_2208_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1192_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1192_in1 = bnn_N_Mux_2_2_3_1_2208_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1192_in1 = Bline_buffer_60_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1192_in1 = s_reg_905;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1192
         assign bnn_Minus_2S_2S_1_1192_out1 = -bnn_Minus_2S_2S_1_1192_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1193
         assign bnn_Add_4Sx2S_5S_1_1193_out1 = {bnn_Add_4Sx2S_4S_1_1175_out1[3], bnn_Add_4Sx2S_4S_1_1175_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1174_out1[1]}}, bnn_N_Mux_2_2_3_1_1174_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_45_mi61 or s_reg_1112 or s_reg_929 or s_reg_991 or bnn_N_Mux_64_2_2_1_1636_out1[44] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1194_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1194_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[44], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1194_in3 = Bline_buffer_45_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1194_in3 = s_reg_991;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1194_in3 = s_reg_929;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1176_out1 or bnn_N_Mux_2_2_3_1_1194_in3)
          begin :bnn_N_Mux_2_2_3_1_1194
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1194_out1 = bnn_Minus_2S_2S_1_1176_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1194_out1 = bnn_N_Mux_2_2_3_1_1194_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1195
         assign bnn_Add_4Sx2S_4S_1_1195_out1 = bnn_Add_4Sx2S_4S_1_1178_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1177_out1[1]}}, bnn_N_Mux_2_2_3_1_1177_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_46_mi61 or s_reg_1112 or s_reg_936 or s_reg_993 or bnn_N_Mux_64_2_2_1_1636_out1[45] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1196_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1196_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1196_in1 = Bline_buffer_46_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1196_in1 = s_reg_993;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1196_in1 = s_reg_936;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1196
         assign bnn_Minus_2S_2S_1_1196_out1 = -bnn_Minus_2S_2S_1_1196_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1179_out1 or bnn_N_Mux_2_2_3_1_1194_in3)
          begin :bnn_N_Mux_2_2_3_1_1197
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1197_out1 = bnn_Minus_2S_2S_1_1179_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1197_out1 = bnn_N_Mux_2_2_3_1_1194_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1198
         assign bnn_Add_4Sx2S_4S_1_1198_out1 = bnn_Add_3Sx3S_4S_1_1181_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1180_out1[1]}}, bnn_N_Mux_2_2_3_1_1180_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1199
         assign bnn_Minus_2S_2S_1_1199_out1 = -bnn_Minus_2S_2S_1_1196_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1182_out1 or bnn_N_Mux_2_2_3_1_1194_in3)
          begin :bnn_N_Mux_2_2_3_1_1200
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1200_out1 = bnn_Minus_2S_2S_1_1182_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1200_out1 = bnn_N_Mux_2_2_3_1_1194_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1201
         assign bnn_Add_3Sx3S_4S_1_1201_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1184_out1[1]}}, bnn_N_Mux_2_2_3_1_1184_out1} + {bnn_Add_2Sx2S_3S_1_1183_out1[2], bnn_Add_2Sx2S_3S_1_1183_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_46_mi61 or s_reg_1112 or s_reg_936 or bnn_N_Mux_64_2_2_1_1636_out1[45] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1202_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1202_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1202_in1 = Bline_buffer_46_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1202_in1 = s_reg_936;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1202
         assign bnn_Minus_2S_2S_4_1202_out1 = -bnn_Minus_2S_2S_4_1202_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1203
         assign bnn_Add_2Sx2S_3S_1_1203_out1 = {bnn_N_Mux_2_2_3_1_1186_out1[1], bnn_N_Mux_2_2_3_1_1186_out1} + {bnn_N_Mux_2_2_3_1_1185_out1[1], bnn_N_Mux_2_2_3_1_1185_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1187_out1 or bnn_N_Mux_2_2_3_1_1188_in3)
          begin :bnn_N_Mux_2_2_3_1_1204
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1204_out1 = bnn_Minus_2S_2S_1_1187_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1204_out1 = bnn_N_Mux_2_2_3_1_1188_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_47_mi61 or s_reg_1112 or s_reg_940 or bnn_N_Mux_64_2_2_1_1636_out1[46] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1205_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1205_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1205_in1 = Bline_buffer_47_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1205_in1 = s_reg_940;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1205
         assign bnn_Minus_2S_2S_4_1205_out1 = -bnn_Minus_2S_2S_4_1205_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1206
         assign bnn_Add_2Sx2S_3S_1_1206_out1 = {bnn_N_Mux_2_2_3_1_1189_out1[1], bnn_N_Mux_2_2_3_1_1189_out1} + {bnn_N_Mux_2_2_3_1_1188_out1[1], bnn_N_Mux_2_2_3_1_1188_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_39_mi61 or s_reg_1112 or s_reg_935 or bnn_N_Mux_2_2_3_1_2190_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1207_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1207_in3 = bnn_N_Mux_2_2_3_1_2190_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1207_in3 = Bline_buffer_39_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1207_in3 = s_reg_935;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1190_out1 or bnn_N_Mux_2_2_3_1_1207_in3)
          begin :bnn_N_Mux_2_2_3_1_1207
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1207_out1 = bnn_Minus_2S_2S_1_1190_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1207_out1 = bnn_N_Mux_2_2_3_1_1207_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_61_mi61 or s_reg_1112 or s_reg_896 or bnn_N_Mux_2_2_3_1_2021_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1208_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1208_in3 = bnn_N_Mux_2_2_3_1_2021_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1208_in3 = Bline_buffer_61_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1208_in3 = s_reg_896;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1191_out1 or bnn_N_Mux_2_2_3_1_1208_in3)
          begin :bnn_N_Mux_2_2_3_1_1208
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1208_out1 = bnn_Minus_2S_2S_1_1191_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1208_out1 = bnn_N_Mux_2_2_3_1_1208_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_60_mi61 or s_reg_1112 or s_reg_905 or bnn_N_Mux_2_2_3_1_2208_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1209_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1209_in3 = bnn_N_Mux_2_2_3_1_2208_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1209_in3 = Bline_buffer_60_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1209_in3 = s_reg_905;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_Minus_2S_2S_1_1192_out1 or bnn_N_Mux_2_2_3_1_1209_in3)
          begin :bnn_N_Mux_2_2_3_1_1209
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1209_out1 = bnn_Minus_2S_2S_1_1192_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1209_out1 = bnn_N_Mux_2_2_3_1_1209_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_62_mi61 or s_reg_1112 or s_reg_906 or bnn_N_Mux_2_2_3_1_2038_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1210_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1210_in1 = bnn_N_Mux_2_2_3_1_2038_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1210_in1 = Bline_buffer_62_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1210_in1 = s_reg_906;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1210
         assign bnn_Minus_2S_2S_1_1210_out1 = -bnn_Minus_2S_2S_1_1210_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1211
         assign bnn_Add_4Sx2S_5S_1_1211_out1 = {bnn_Add_4Sx2S_4S_1_1195_out1[3], bnn_Add_4Sx2S_4S_1_1195_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1194_out1[1]}}, bnn_N_Mux_2_2_3_1_1194_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_46_mi61 or s_reg_1112 or s_reg_936 or s_reg_993 or bnn_N_Mux_64_2_2_1_1636_out1[45] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1212_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1212_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1212_in3 = Bline_buffer_46_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1212_in3 = s_reg_993;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1212_in3 = s_reg_936;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1196_out1 or bnn_N_Mux_2_2_3_1_1212_in3)
          begin :bnn_N_Mux_2_2_3_1_1212
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1212_out1 = bnn_Minus_2S_2S_1_1196_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1212_out1 = bnn_N_Mux_2_2_3_1_1212_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1213
         assign bnn_Add_4Sx2S_4S_1_1213_out1 = bnn_Add_4Sx2S_4S_1_1198_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1197_out1[1]}}, bnn_N_Mux_2_2_3_1_1197_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_47_mi61 or s_reg_1112 or s_reg_940 or s_reg_995 or bnn_N_Mux_64_2_2_1_1636_out1[46] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1214_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1214_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1214_in1 = Bline_buffer_47_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1214_in1 = s_reg_995;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1214_in1 = s_reg_940;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1214
         assign bnn_Minus_2S_2S_1_1214_out1 = -bnn_Minus_2S_2S_1_1214_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1199_out1 or bnn_N_Mux_2_2_3_1_1212_in3)
          begin :bnn_N_Mux_2_2_3_1_1215
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1215_out1 = bnn_Minus_2S_2S_1_1199_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1215_out1 = bnn_N_Mux_2_2_3_1_1212_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1216
         assign bnn_Add_4Sx2S_4S_1_1216_out1 = bnn_Add_3Sx3S_4S_1_1201_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1200_out1[1]}}, bnn_N_Mux_2_2_3_1_1200_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1217
         assign bnn_Minus_2S_2S_4_1217_out1 = -bnn_Minus_2S_2S_4_1205_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_46_mi61 or s_reg_1112 or s_reg_936 or bnn_N_Mux_64_2_2_1_1636_out1[45] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1218_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1218_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1218_in3 = Bline_buffer_46_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1218_in3 = s_reg_936;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1202_out1 or bnn_N_Mux_2_2_3_4_1218_in3)
          begin :bnn_N_Mux_2_2_3_4_1218
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1218_out1 = bnn_Minus_2S_2S_4_1202_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1218_out1 = bnn_N_Mux_2_2_3_4_1218_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1219
         assign bnn_Add_3Sx3S_4S_1_1219_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1204_out1[1]}}, bnn_N_Mux_2_2_3_1_1204_out1} + {bnn_Add_2Sx2S_3S_1_1203_out1[2], bnn_Add_2Sx2S_3S_1_1203_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1220
         assign bnn_Minus_2S_2S_1_1220_out1 = -bnn_Minus_2S_2S_1_1210_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1221
         assign bnn_Minus_2S_2S_1_1221_out1 = -bnn_Minus_2S_2S_1_1191_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_48_mi61 or s_reg_1112 or s_reg_945 or bnn_N_Mux_64_2_2_1_1636_out1[47] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1222_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1222_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[47], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1222_in1 = Bline_buffer_48_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1222_in1 = s_reg_945;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1222
         assign bnn_Minus_2S_2S_4_1222_out1 = -bnn_Minus_2S_2S_4_1222_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_47_mi61 or s_reg_1112 or s_reg_940 or bnn_N_Mux_64_2_2_1_1636_out1[46] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1223_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1223_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1223_in3 = Bline_buffer_47_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1223_in3 = s_reg_940;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1205_out1 or bnn_N_Mux_2_2_3_4_1223_in3)
          begin :bnn_N_Mux_2_2_3_4_1223
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1223_out1 = bnn_Minus_2S_2S_4_1205_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1223_out1 = bnn_N_Mux_2_2_3_4_1223_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1224
         assign bnn_Add_3Sx3S_4S_1_1224_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1207_out1[1]}}, bnn_N_Mux_2_2_3_1_1207_out1} + {bnn_Add_2Sx2S_3S_1_1206_out1[2], bnn_Add_2Sx2S_3S_1_1206_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_70_mi61 or s_reg_1112 or s_reg_948 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1640_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_1225_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1225_in1 = bnn_N_Mux_3_2_6_4_1640_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_1225_in1 = Bline_buffer_70_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1225_in1 = s_reg_948;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1225
         assign bnn_Minus_2S_2S_4_1225_out1 = -bnn_Minus_2S_2S_4_1225_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1226
         assign bnn_Add_2Sx2S_3S_1_1226_out1 = {bnn_N_Mux_2_2_3_1_1209_out1[1], bnn_N_Mux_2_2_3_1_1209_out1} + {bnn_N_Mux_2_2_3_1_1208_out1[1], bnn_N_Mux_2_2_3_1_1208_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_62_mi61 or s_reg_1112 or s_reg_906 or bnn_N_Mux_2_2_3_1_2038_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1227_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1227_in3 = bnn_N_Mux_2_2_3_1_2038_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1227_in3 = Bline_buffer_62_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1227_in3 = s_reg_906;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1210_out1 or bnn_N_Mux_2_2_3_1_1227_in3)
          begin :bnn_N_Mux_2_2_3_1_1227
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1227_out1 = bnn_Minus_2S_2S_1_1210_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1227_out1 = bnn_N_Mux_2_2_3_1_1227_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1228
         assign bnn_Add_4Sx2S_5S_1_1228_out1 = {bnn_Add_4Sx2S_4S_1_1213_out1[3], bnn_Add_4Sx2S_4S_1_1213_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1212_out1[1]}}, bnn_N_Mux_2_2_3_1_1212_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_47_mi61 or s_reg_1112 or s_reg_940 or s_reg_995 or bnn_N_Mux_64_2_2_1_1636_out1[46] or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1229_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1229_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1229_in3 = Bline_buffer_47_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1229_in3 = s_reg_995;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1229_in3 = s_reg_940;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_1214_out1 or bnn_N_Mux_2_2_3_1_1229_in3)
          begin :bnn_N_Mux_2_2_3_1_1229
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_1229_out1 = bnn_Minus_2S_2S_1_1214_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1229_out1 = bnn_N_Mux_2_2_3_1_1229_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1230
         assign bnn_Add_4Sx2S_4S_1_1230_out1 = bnn_Add_4Sx2S_4S_1_1216_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1215_out1[1]}}, bnn_N_Mux_2_2_3_1_1215_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1231
         assign bnn_Minus_2S_2S_4_1231_out1 = -bnn_Minus_2S_2S_4_1222_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1217_out1 or bnn_N_Mux_2_2_3_4_1223_in3)
          begin :bnn_N_Mux_2_2_3_4_1232
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1232_out1 = bnn_Minus_2S_2S_4_1217_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1232_out1 = bnn_N_Mux_2_2_3_4_1223_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1233
         assign bnn_Add_4Sx2S_4S_1_1233_out1 = bnn_Add_3Sx3S_4S_1_1219_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1218_out1[1]}}, bnn_N_Mux_2_2_3_4_1218_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1220_out1 or bnn_N_Mux_2_2_3_1_1227_in3)
          begin :bnn_N_Mux_2_2_3_1_1234
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1234_out1 = bnn_Minus_2S_2S_1_1220_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1234_out1 = bnn_N_Mux_2_2_3_1_1227_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1208_in3 or bnn_Minus_2S_2S_1_1221_out1)
          begin :bnn_N_Mux_2_2_3_1_1235
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1235_out1 = bnn_Minus_2S_2S_1_1221_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1235_out1 = bnn_N_Mux_2_2_3_1_1208_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_63_mi61 or s_reg_1112 or s_reg_915 or bnn_N_Mux_2_2_3_1_2055_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1236_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1236_in1 = bnn_N_Mux_2_2_3_1_2055_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1236_in1 = Bline_buffer_63_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1236_in1 = s_reg_915;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1236
         assign bnn_Minus_2S_2S_1_1236_out1 = -bnn_Minus_2S_2S_1_1236_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1237
         assign bnn_Minus_2S_2S_1_1237_out1 = -bnn_Minus_2S_2S_1_1236_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1238
         assign bnn_Minus_2S_2S_1_1238_out1 = -bnn_Minus_2S_2S_1_1210_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_49_mi61 or s_reg_1112 or s_reg_952 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_1_1639_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_1239_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1239_in1 = bnn_N_Mux_3_2_6_1_1639_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_1239_in1 = Bline_buffer_49_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1239_in1 = s_reg_952;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1239
         assign bnn_Minus_2S_2S_4_1239_out1 = -bnn_Minus_2S_2S_4_1239_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_48_mi61 or s_reg_1112 or s_reg_945 or bnn_N_Mux_64_2_2_1_1636_out1[47] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1240_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1240_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[47], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1240_in3 = Bline_buffer_48_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1240_in3 = s_reg_945;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1222_out1 or bnn_N_Mux_2_2_3_4_1240_in3)
          begin :bnn_N_Mux_2_2_3_4_1240
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1240_out1 = bnn_Minus_2S_2S_4_1222_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1240_out1 = bnn_N_Mux_2_2_3_4_1240_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1241
         assign bnn_Add_4Sx2S_4S_1_1241_out1 = bnn_Add_3Sx3S_4S_1_1224_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1223_out1[1]}}, bnn_N_Mux_2_2_3_4_1223_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_71_mi61 or s_reg_1112 or s_reg_954 or bnn_N_Mux_64_2_2_1_1636_out1[48] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1242_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1242_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[48], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1242_in1 = Bline_buffer_71_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1242_in1 = s_reg_954;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1242
         assign bnn_Minus_2S_2S_4_1242_out1 = -bnn_Minus_2S_2S_4_1242_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_70_mi61 or s_reg_1112 or s_reg_948 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_1640_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_1243_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1243_in3 = bnn_N_Mux_3_2_6_4_1640_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1243_in3 = Bline_buffer_70_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1243_in3 = s_reg_948;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1225_out1 or bnn_N_Mux_2_2_3_4_1243_in3)
          begin :bnn_N_Mux_2_2_3_4_1243
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1243_out1 = bnn_Minus_2S_2S_4_1225_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1243_out1 = bnn_N_Mux_2_2_3_4_1243_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1244
         assign bnn_Add_3Sx3S_4S_1_1244_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1227_out1[1]}}, bnn_N_Mux_2_2_3_1_1227_out1} + {bnn_Add_2Sx2S_3S_1_1226_out1[2], bnn_Add_2Sx2S_3S_1_1226_out1};

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1245
         assign bnn_Add_4Sx2S_5S_1_1245_out1 = {bnn_Add_4Sx2S_4S_1_1230_out1[3], bnn_Add_4Sx2S_4S_1_1230_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_1229_out1[1]}}, bnn_N_Mux_2_2_3_1_1229_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1231_out1 or bnn_N_Mux_2_2_3_4_1240_in3)
          begin :bnn_N_Mux_2_2_3_4_1246
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1246_out1 = bnn_Minus_2S_2S_4_1231_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1246_out1 = bnn_N_Mux_2_2_3_4_1240_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1247
         assign bnn_Add_4Sx2S_4S_1_1247_out1 = bnn_Add_4Sx2S_4S_1_1233_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1232_out1[1]}}, bnn_N_Mux_2_2_3_4_1232_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1248
         assign bnn_Minus_2S_2S_4_1248_out1 = -bnn_Minus_2S_2S_4_1242_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1249
         assign bnn_Add_2Sx2S_3S_1_1249_out1 = {bnn_N_Mux_2_2_3_1_1235_out1[1], bnn_N_Mux_2_2_3_1_1235_out1} + {bnn_N_Mux_2_2_3_1_1234_out1[1], bnn_N_Mux_2_2_3_1_1234_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_63_mi61 or s_reg_1112 or s_reg_915 or bnn_N_Mux_2_2_3_1_2055_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1250_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1250_in3 = bnn_N_Mux_2_2_3_1_2055_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1250_in3 = Bline_buffer_63_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1250_in3 = s_reg_915;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_1236_out1 or bnn_N_Mux_2_2_3_1_1250_in3)
          begin :bnn_N_Mux_2_2_3_1_1250
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1250_out1 = bnn_Minus_2S_2S_1_1236_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1250_out1 = bnn_N_Mux_2_2_3_1_1250_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1237_out1 or bnn_N_Mux_2_2_3_1_1250_in3)
          begin :bnn_N_Mux_2_2_3_1_1251
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1251_out1 = bnn_Minus_2S_2S_1_1237_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1251_out1 = bnn_N_Mux_2_2_3_1_1250_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1227_in3 or bnn_Minus_2S_2S_1_1238_out1)
          begin :bnn_N_Mux_2_2_3_1_1252
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1252_out1 = bnn_Minus_2S_2S_1_1238_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1252_out1 = bnn_N_Mux_2_2_3_1_1227_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_64_mi61 or s_reg_1112 or s_reg_923 or bnn_N_Mux_2_2_3_1_2072_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1253_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1253_in1 = bnn_N_Mux_2_2_3_1_2072_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1253_in1 = Bline_buffer_64_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1253_in1 = s_reg_923;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1253
         assign bnn_Minus_2S_2S_4_1253_out1 = -bnn_Minus_2S_2S_4_1253_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1254
         assign bnn_Minus_2S_2S_4_1254_out1 = -bnn_Minus_2S_2S_4_1253_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1255
         assign bnn_Minus_2S_2S_4_1255_out1 = -bnn_Minus_2S_2S_1_1236_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_49_mi61 or s_reg_1112 or s_reg_952 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_1_1639_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_1256_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1256_in3 = bnn_N_Mux_3_2_6_1_1639_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1256_in3 = Bline_buffer_49_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1256_in3 = s_reg_952;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1239_out1 or bnn_N_Mux_2_2_3_4_1256_in3)
          begin :bnn_N_Mux_2_2_3_4_1256
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1256_out1 = bnn_Minus_2S_2S_4_1239_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1256_out1 = bnn_N_Mux_2_2_3_4_1256_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1257
         assign bnn_Add_4Sx2S_4S_1_1257_out1 = bnn_Add_4Sx2S_4S_1_1241_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1240_out1[1]}}, bnn_N_Mux_2_2_3_4_1240_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_72_mi61 or s_reg_1112 or s_reg_958 or bnn_N_Mux_64_2_2_1_1636_out1[49] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1258_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1258_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[49], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1258_in1 = Bline_buffer_72_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1258_in1 = s_reg_958;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1258
         assign bnn_Minus_2S_2S_4_1258_out1 = -bnn_Minus_2S_2S_4_1258_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_71_mi61 or s_reg_1112 or s_reg_954 or bnn_N_Mux_64_2_2_1_1636_out1[48] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1259_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1259_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[48], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1259_in3 = Bline_buffer_71_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1259_in3 = s_reg_954;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1242_out1 or bnn_N_Mux_2_2_3_4_1259_in3)
          begin :bnn_N_Mux_2_2_3_4_1259
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1259_out1 = bnn_Minus_2S_2S_4_1242_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1259_out1 = bnn_N_Mux_2_2_3_4_1259_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1260
         assign bnn_Add_4Sx2S_4S_1_1260_out1 = bnn_Add_3Sx3S_4S_1_1244_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1243_out1[1]}}, bnn_N_Mux_2_2_3_4_1243_out1};

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1261
         assign bnn_Add_4Sx2S_5S_1_1261_out1 = {bnn_Add_4Sx2S_4S_1_1247_out1[3], bnn_Add_4Sx2S_4S_1_1247_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1246_out1[1]}}, bnn_N_Mux_2_2_3_4_1246_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1248_out1 or bnn_N_Mux_2_2_3_4_1259_in3)
          begin :bnn_N_Mux_2_2_3_4_1262
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1262_out1 = bnn_Minus_2S_2S_4_1248_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1262_out1 = bnn_N_Mux_2_2_3_4_1259_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1263
         assign bnn_Add_3Sx3S_4S_1_1263_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1250_out1[1]}}, bnn_N_Mux_2_2_3_1_1250_out1} + {bnn_Add_2Sx2S_3S_1_1249_out1[2], bnn_Add_2Sx2S_3S_1_1249_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1264
         assign bnn_Add_2Sx2S_3S_1_1264_out1 = {bnn_N_Mux_2_2_3_1_1252_out1[1], bnn_N_Mux_2_2_3_1_1252_out1} + {bnn_N_Mux_2_2_3_1_1251_out1[1], bnn_N_Mux_2_2_3_1_1251_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_64_mi61 or s_reg_1112 or s_reg_923 or bnn_N_Mux_2_2_3_1_2072_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1265_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1265_in3 = bnn_N_Mux_2_2_3_1_2072_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1265_in3 = Bline_buffer_64_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1265_in3 = s_reg_923;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_Minus_2S_2S_4_1253_out1 or bnn_N_Mux_2_2_3_4_1265_in3)
          begin :bnn_N_Mux_2_2_3_4_1265
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_1265_out1 = bnn_Minus_2S_2S_4_1253_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1265_out1 = bnn_N_Mux_2_2_3_4_1265_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_Minus_2S_2S_4_1254_out1 or bnn_N_Mux_2_2_3_4_1265_in3)
          begin :bnn_N_Mux_2_2_3_4_1266
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_1266_out1 = bnn_Minus_2S_2S_4_1254_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1266_out1 = bnn_N_Mux_2_2_3_4_1265_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1250_in3 or bnn_Minus_2S_2S_4_1255_out1)
          begin :bnn_N_Mux_2_2_3_4_1267
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1267_out1 = bnn_Minus_2S_2S_4_1255_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1267_out1 = bnn_N_Mux_2_2_3_1_1250_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1268
         assign bnn_Minus_2S_2S_4_1268_out1 = -bnn_Minus_2S_2S_4_1253_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1269
         assign bnn_Add_4Sx2S_5S_1_1269_out1 = {bnn_Add_4Sx2S_4S_1_1257_out1[3], bnn_Add_4Sx2S_4S_1_1257_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1256_out1[1]}}, bnn_N_Mux_2_2_3_4_1256_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_72_mi61 or s_reg_1112 or s_reg_958 or bnn_N_Mux_64_2_2_1_1636_out1[49] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1270_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1270_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[49], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1270_in3 = Bline_buffer_72_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1270_in3 = s_reg_958;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1258_out1 or bnn_N_Mux_2_2_3_4_1270_in3)
          begin :bnn_N_Mux_2_2_3_4_1270
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1270_out1 = bnn_Minus_2S_2S_4_1258_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1270_out1 = bnn_N_Mux_2_2_3_4_1270_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1271
         assign bnn_Add_4Sx2S_4S_1_1271_out1 = bnn_Add_4Sx2S_4S_1_1260_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1259_out1[1]}}, bnn_N_Mux_2_2_3_4_1259_out1};

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1272
         assign bnn_Add_4Sx2S_4S_1_1272_out1 = bnn_Add_3Sx3S_4S_1_1263_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1262_out1[1]}}, bnn_N_Mux_2_2_3_4_1262_out1};

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1273
         assign bnn_Add_3Sx3S_4S_1_1273_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1265_out1[1]}}, bnn_N_Mux_2_2_3_4_1265_out1} + {bnn_Add_2Sx2S_3S_1_1264_out1[2], bnn_Add_2Sx2S_3S_1_1264_out1};

         // resource: bnn_Add_2Sx2S_3S_4  instance: bnn_Add_2Sx2S_3S_4_1274
         assign bnn_Add_2Sx2S_3S_4_1274_out1 = {bnn_N_Mux_2_2_3_4_1267_out1[1], bnn_N_Mux_2_2_3_4_1267_out1} + {bnn_N_Mux_2_2_3_4_1266_out1[1], bnn_N_Mux_2_2_3_4_1266_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1275
         assign bnn_Minus_2S_2S_4_1275_out1 = -bnn_Minus_2S_2S_4_1258_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1276
         assign bnn_Minus_2S_2S_4_1276_out1 = -bnn_Minus_2S_2S_4_1258_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_N_Mux_2_2_3_4_1270_in3 or bnn_Minus_2S_2S_4_1275_out1)
          begin :bnn_N_Mux_2_2_3_4_1277
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1277_out1 = bnn_Minus_2S_2S_4_1275_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1277_out1 = bnn_N_Mux_2_2_3_4_1270_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_N_Mux_2_2_3_4_1270_in3 or bnn_Minus_2S_2S_4_1276_out1)
          begin :bnn_N_Mux_2_2_3_4_1278
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1278_out1 = bnn_Minus_2S_2S_4_1276_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1278_out1 = bnn_N_Mux_2_2_3_4_1270_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_4_1265_in3 or bnn_Minus_2S_2S_4_1268_out1)
          begin :bnn_N_Mux_2_2_3_4_1279
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1279_out1 = bnn_Minus_2S_2S_4_1268_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1279_out1 = bnn_N_Mux_2_2_3_4_1265_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1280
         assign bnn_Add_4Sx2S_5S_1_1280_out1 = {bnn_Add_4Sx2S_4S_1_1271_out1[3], bnn_Add_4Sx2S_4S_1_1271_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1270_out1[1]}}, bnn_N_Mux_2_2_3_4_1270_out1};

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1281
         assign bnn_Add_4Sx2S_4S_1_1281_out1 = bnn_Add_4Sx2S_4S_1_1272_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1277_out1[1]}}, bnn_N_Mux_2_2_3_4_1277_out1};

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1282
         assign bnn_Add_4Sx3S_4S_1_1282_out1 = bnn_Add_3Sx3S_4S_1_1273_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1278_out1[1]}}, bnn_N_Mux_2_2_3_4_1278_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_68_mi61 or s_reg_1112 or s_reg_947 or bnn_N_Mux_2_2_3_1_2140_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1283_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1283_in1 = bnn_N_Mux_2_2_3_1_2140_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1283_in1 = Bline_buffer_68_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1283_in1 = s_reg_947;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1283
         assign bnn_Minus_2S_2S_4_1283_out1 = -bnn_Minus_2S_2S_4_1283_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_67_mi61 or s_reg_1112 or s_reg_942 or bnn_N_Mux_2_2_3_1_2123_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1284_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1284_in1 = bnn_N_Mux_2_2_3_1_2123_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1284_in1 = Bline_buffer_67_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1284_in1 = s_reg_942;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1284
         assign bnn_Minus_2S_2S_4_1284_out1 = -bnn_Minus_2S_2S_4_1284_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_68_mi61 or s_reg_1112 or s_reg_947 or bnn_N_Mux_2_2_3_1_2140_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1285_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1285_in3 = bnn_N_Mux_2_2_3_1_2140_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1285_in3 = Bline_buffer_68_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1285_in3 = s_reg_947;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_Minus_2S_2S_4_1283_out1 or bnn_N_Mux_2_2_3_4_1285_in3)
          begin :bnn_N_Mux_2_2_3_4_1285
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_1285_out1 = bnn_Minus_2S_2S_4_1283_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1285_out1 = bnn_N_Mux_2_2_3_4_1285_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_67_mi61 or s_reg_1112 or s_reg_942 or bnn_N_Mux_2_2_3_1_2123_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1286_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1286_in3 = bnn_N_Mux_2_2_3_1_2123_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1286_in3 = Bline_buffer_67_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1286_in3 = s_reg_942;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_Minus_2S_2S_4_1284_out1 or bnn_N_Mux_2_2_3_4_1286_in3)
          begin :bnn_N_Mux_2_2_3_4_1286
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1286_out1 = bnn_Minus_2S_2S_4_1284_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1286_out1 = bnn_N_Mux_2_2_3_4_1286_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_69_mi61 or s_reg_1112 or s_reg_911 or s_reg_971 or bnn_N_Mux_2_2_3_1_3184_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1287_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1287_in1 = bnn_N_Mux_2_2_3_1_3184_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1287_in1 = Bline_buffer_69_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1287_in1 = s_reg_971;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1287_in1 = s_reg_911;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1287
         assign bnn_Minus_2S_2S_1_1287_out1 = -bnn_Minus_2S_2S_1_1287_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_91_mi61 or s_reg_1112 or s_reg_927 or bnn_N_Mux_2_2_3_1_3215_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1288_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1288_in1 = bnn_N_Mux_2_2_3_1_3215_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1288_in1 = Bline_buffer_91_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1288_in1 = s_reg_927;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1288
         assign bnn_Minus_2S_2S_1_1288_out1 = -bnn_Minus_2S_2S_1_1288_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_90_mi61 or s_reg_1112 or s_reg_946 or bnn_N_Mux_2_2_3_1_3337_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1289_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1289_in1 = bnn_N_Mux_2_2_3_1_3337_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1289_in1 = Bline_buffer_90_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1289_in1 = s_reg_946;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1289
         assign bnn_Minus_2S_2S_1_1289_out1 = -bnn_Minus_2S_2S_1_1289_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_77_mi61 or s_reg_1112 or s_reg_873 or s_reg_994 or bnn_N_Mux_2_2_3_1_3093_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1290_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1290_in1 = bnn_N_Mux_2_2_3_1_3093_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1290_in1 = Bline_buffer_77_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1290_in1 = s_reg_994;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1290_in1 = s_reg_873;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1290
         assign bnn_Minus_2S_2S_1_1290_out1 = -bnn_Minus_2S_2S_1_1290_in1;

         // resource: bnn_Add_2Sx2S_3S_4  instance: bnn_Add_2Sx2S_3S_4_1291
         assign bnn_Add_2Sx2S_3S_4_1291_out1 = {bnn_N_Mux_2_2_3_4_1286_out1[1], bnn_N_Mux_2_2_3_4_1286_out1} + {bnn_N_Mux_2_2_3_4_1285_out1[1], bnn_N_Mux_2_2_3_4_1285_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_69_mi61 or s_reg_1112 or s_reg_911 or bnn_N_Mux_2_2_3_1_3184_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1292_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1292_in3 = bnn_N_Mux_2_2_3_1_3184_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1292_in3 = Bline_buffer_69_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1292_in3 = s_reg_911;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_916 or s_reg_951 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1292_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1292_ctrl1 = s_reg_951;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1292_ctrl1 = s_reg_916;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1292_ctrl1 = s_reg_951;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Minus_2S_2S_1_1287_out1 or bnn_N_Mux_2_2_3_4_1292_in3 or bnn_N_Mux_2_2_3_4_1292_ctrl1)
          begin :bnn_N_Mux_2_2_3_4_1292
            if (bnn_N_Mux_2_2_3_4_1292_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1292_out1 = bnn_Minus_2S_2S_1_1287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1292_out1 = bnn_N_Mux_2_2_3_4_1292_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_91_mi61 or s_reg_1112 or s_reg_927 or bnn_N_Mux_2_2_3_1_3215_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1293_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1293_in3 = bnn_N_Mux_2_2_3_1_3215_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1293_in3 = Bline_buffer_91_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1293_in3 = s_reg_927;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_907 or s_reg_957 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1293_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1293_ctrl1 = s_reg_957;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1293_ctrl1 = s_reg_907;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1293_ctrl1 = s_reg_957;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1288_out1 or bnn_N_Mux_2_2_3_1_1293_in3 or bnn_N_Mux_2_2_3_1_1293_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1293
            if (bnn_N_Mux_2_2_3_1_1293_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1293_out1 = bnn_Minus_2S_2S_1_1288_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1293_out1 = bnn_N_Mux_2_2_3_1_1293_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_90_mi61 or s_reg_1112 or s_reg_946 or bnn_N_Mux_2_2_3_1_3337_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1294_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1294_in3 = bnn_N_Mux_2_2_3_1_3337_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1294_in3 = Bline_buffer_90_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1294_in3 = s_reg_946;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_908 or s_reg_957 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1294_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1294_ctrl1 = s_reg_957;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1294_ctrl1 = s_reg_908;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1294_ctrl1 = s_reg_957;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1289_out1 or bnn_N_Mux_2_2_3_1_1294_in3 or bnn_N_Mux_2_2_3_1_1294_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1294
            if (bnn_N_Mux_2_2_3_1_1294_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1294_out1 = bnn_Minus_2S_2S_1_1289_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1294_out1 = bnn_N_Mux_2_2_3_1_1294_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_92_mi61 or s_reg_1112 or s_reg_941 or s_reg_962 or bnn_N_Mux_2_2_3_1_3322_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1295_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1295_in1 = bnn_N_Mux_2_2_3_1_3322_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1295_in1 = Bline_buffer_92_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1295_in1 = s_reg_962;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1295_in1 = s_reg_941;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1295
         assign bnn_Minus_2S_2S_1_1295_out1 = -bnn_Minus_2S_2S_1_1295_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_78_mi61 or s_reg_1112 or s_reg_878 or s_reg_996 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1296_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1296_in1 = bnn_N_Mux_2_2_3_1_3114_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1296_in1 = Bline_buffer_78_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1296_in1 = s_reg_996;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1296_in1 = s_reg_878;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1296
         assign bnn_Minus_2S_2S_1_1296_out1 = -bnn_Minus_2S_2S_1_1296_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(Bline_buffer_77_mi61 or s_reg_924 or bnn_Minus_2S_2S_1_1290_out1)
          begin :bnn_N_Mux_2_2_3_4_1297
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1297_out1 = bnn_Minus_2S_2S_1_1290_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1297_out1 = Bline_buffer_77_mi61;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1298
         assign bnn_Add_3Sx3S_4S_4_1298_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1292_out1[1]}}, bnn_N_Mux_2_2_3_4_1292_out1} + {bnn_Add_2Sx2S_3S_4_1291_out1[2], bnn_Add_2Sx2S_3S_4_1291_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_100_mi61 or s_reg_1112 or s_reg_886[1:0] or s_reg_976 or bnn_N_Mux_2_2_3_1_3216_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1299_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1299_in1 = bnn_N_Mux_2_2_3_1_3216_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1299_in1 = Bline_buffer_100_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1299_in1 = s_reg_976;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1299_in1 = s_reg_886[1:0];
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1299
         assign bnn_Minus_2S_2S_1_1299_out1 = -bnn_Minus_2S_2S_1_1299_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1300
         assign bnn_Add_2Sx2S_3S_1_1300_out1 = {bnn_N_Mux_2_2_3_1_1294_out1[1], bnn_N_Mux_2_2_3_1_1294_out1} + {bnn_N_Mux_2_2_3_1_1293_out1[1], bnn_N_Mux_2_2_3_1_1293_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_92_mi61 or s_reg_1112 or s_reg_941 or bnn_N_Mux_2_2_3_1_3322_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1301_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1301_in3 = bnn_N_Mux_2_2_3_1_3322_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1301_in3 = Bline_buffer_92_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1301_in3 = s_reg_941;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_4_1292_ctrl1 or bnn_Minus_2S_2S_1_1295_out1 or bnn_N_Mux_2_2_3_1_1301_in3)
          begin :bnn_N_Mux_2_2_3_1_1301
            if (bnn_N_Mux_2_2_3_4_1292_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1301_out1 = bnn_Minus_2S_2S_1_1295_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1301_out1 = bnn_N_Mux_2_2_3_1_1301_in3;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_79_mi61 or s_reg_1112 or s_reg_872 or s_reg_992 or bnn_N_Mux_2_2_3_1_3071_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1302_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1302_in1 = bnn_N_Mux_2_2_3_1_3071_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1302_in1 = Bline_buffer_79_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1302_in1 = s_reg_992;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1302_in1 = s_reg_872;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1302
         assign bnn_Minus_2S_2S_1_1302_out1 = -bnn_Minus_2S_2S_1_1302_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(Bline_buffer_78_mi61 or s_reg_932 or bnn_Minus_2S_2S_1_1296_out1)
          begin :bnn_N_Mux_2_2_3_4_1303
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1303_out1 = bnn_Minus_2S_2S_1_1296_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1303_out1 = Bline_buffer_78_mi61;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1304
         assign bnn_Add_4Sx3S_4S_1_1304_out1 = bnn_Add_3Sx3S_4S_4_1298_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1297_out1[1]}}, bnn_N_Mux_2_2_3_4_1297_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_101_mi61 or s_reg_1112 or s_reg_878 or s_reg_998 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1305_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1305_in1 = bnn_N_Mux_2_2_3_1_3114_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1305_in1 = Bline_buffer_101_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1305_in1 = s_reg_998;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1305_in1 = s_reg_878;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1305
         assign bnn_Minus_2S_2S_1_1305_out1 = -bnn_Minus_2S_2S_1_1305_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_100_mi61 or s_reg_1112 or s_reg_886[1:0] or s_reg_976 or bnn_N_Mux_2_2_3_1_3216_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1306_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1306_in3 = bnn_N_Mux_2_2_3_1_3216_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1306_in3 = Bline_buffer_100_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1306_in3 = s_reg_976;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1306_in3 = s_reg_886[1:0];
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_924 or s_reg_944 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1306_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1306_ctrl1 = s_reg_944;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1306_ctrl1 = s_reg_924;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1306_ctrl1 = s_reg_944;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1299_out1 or bnn_N_Mux_2_2_3_1_1306_in3 or bnn_N_Mux_2_2_3_1_1306_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1306
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1306_out1 = bnn_Minus_2S_2S_1_1299_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1306_out1 = bnn_N_Mux_2_2_3_1_1306_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1307
         assign bnn_Add_3Sx3S_4S_1_1307_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1301_out1[1]}}, bnn_N_Mux_2_2_3_1_1301_out1} + {bnn_Add_2Sx2S_3S_1_1300_out1[2], bnn_Add_2Sx2S_3S_1_1300_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_79_mi61 or s_reg_1112 or s_reg_872 or bnn_N_Mux_2_2_3_1_3071_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1308_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1308_in3 = bnn_N_Mux_2_2_3_1_3071_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1308_in3 = Bline_buffer_79_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1308_in3 = s_reg_872;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_939 or s_reg_951 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1308_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1308_ctrl1 = s_reg_951;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1308_ctrl1 = s_reg_939;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1308_ctrl1 = s_reg_951;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Minus_2S_2S_1_1302_out1 or bnn_N_Mux_2_2_3_4_1308_in3 or bnn_N_Mux_2_2_3_4_1308_ctrl1)
          begin :bnn_N_Mux_2_2_3_4_1308
            if (bnn_N_Mux_2_2_3_4_1308_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1308_out1 = bnn_Minus_2S_2S_1_1302_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1308_out1 = bnn_N_Mux_2_2_3_4_1308_in3;
            end
         end

         // resource: mux_4bx2i
         always @(s_reg_1112 or bnn_Add_4Sx3S_4S_1_1017_out1 or bnn_Add_4Sx3S_4S_1_1304_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_4Sx2S_5S_4_1309_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_4Sx2S_5S_4_1309_in2 = bnn_Add_4Sx3S_4S_1_1017_out1;
               end
               else begin
                  bnn_Add_4Sx2S_5S_4_1309_in2 = bnn_Add_4Sx3S_4S_1_1304_out1;
               end
            end
            else begin
               bnn_Add_4Sx2S_5S_4_1309_in2 = bnn_Add_4Sx3S_4S_1_1017_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_4_1303_out1 or bnn_N_Mux_2_2_3_4_1486_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_4Sx2S_5S_4_1309_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_4Sx2S_5S_4_1309_in1 = bnn_N_Mux_2_2_3_4_1486_out1;
               end
               else begin
                  bnn_Add_4Sx2S_5S_4_1309_in1 = bnn_N_Mux_2_2_3_4_1303_out1;
               end
            end
            else begin
               bnn_Add_4Sx2S_5S_4_1309_in1 = bnn_N_Mux_2_2_3_4_1486_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1309
         assign bnn_Add_4Sx2S_5S_4_1309_out1 = {bnn_Add_4Sx2S_5S_4_1309_in2[3], bnn_Add_4Sx2S_5S_4_1309_in2} + {{ 3 {bnn_Add_4Sx2S_5S_4_1309_in1[1]}}, bnn_Add_4Sx2S_5S_4_1309_in1};

         // resource: mux_2bx4i
         always @(Bline_buffer_102_mi61 or s_reg_1112 or s_reg_895 or s_reg_982 or bnn_N_Mux_2_2_3_1_3229_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1310_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1310_in1 = bnn_N_Mux_2_2_3_1_3229_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1310_in1 = Bline_buffer_102_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1310_in1 = s_reg_982;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1310_in1 = s_reg_895;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1310
         assign bnn_Minus_2S_2S_1_1310_out1 = -bnn_Minus_2S_2S_1_1310_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_101_mi61 or s_reg_1112 or s_reg_878 or s_reg_998 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1311_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1311_in3 = bnn_N_Mux_2_2_3_1_3114_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1311_in3 = Bline_buffer_101_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1311_in3 = s_reg_998;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1311_in3 = s_reg_878;
               end
               
            endcase

         end

         // resource: mux_1bx3i
         always @(s_reg_1112 or s_reg_932 or s_reg_944 or s_reg_951 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1311_ctrl1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1311_ctrl1 = s_reg_944;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1311_ctrl1 = s_reg_932;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1311_ctrl1 = s_reg_951;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1311_ctrl1 = s_reg_944;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1305_out1 or bnn_N_Mux_2_2_3_1_1311_in3 or bnn_N_Mux_2_2_3_1_1311_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1311
            if (bnn_N_Mux_2_2_3_1_1311_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1311_out1 = bnn_Minus_2S_2S_1_1305_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1311_out1 = bnn_N_Mux_2_2_3_1_1311_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1312
         assign bnn_Add_4Sx2S_4S_1_1312_out1 = bnn_Add_3Sx3S_4S_1_1307_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1306_out1[1]}}, bnn_N_Mux_2_2_3_1_1306_out1};

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_4_1309_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_4_1313_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_4_1313_in2 = bnn_Add_4Sx2S_5S_4_1309_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_4_1313_in2 = {bnn_Add_4Sx2S_5S_4_1309_out1[3], bnn_Add_4Sx2S_5S_4_1309_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_4_1313_in2 = bnn_Add_4Sx2S_5S_4_1309_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1313
         assign bnn_Add_5Sx4S_6S_4_1313_out1 = {bnn_Add_5Sx4S_6S_4_1313_in2[4], bnn_Add_5Sx4S_6S_4_1313_in2} + {{ 4 {bnn_N_Mux_2_2_3_4_1308_out1[1]}}, bnn_N_Mux_2_2_3_4_1308_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_102_mi61 or s_reg_1112 or s_reg_884 or bnn_N_Mux_2_2_3_1_3133_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1314_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1314_in3 = bnn_N_Mux_2_2_3_1_3133_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1314_in3 = Bline_buffer_102_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1314_in3 = s_reg_884;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_Minus_2S_2S_1_1310_out1 or bnn_Minus_2S_2S_1_1440_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1314_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1314_in2 = bnn_Minus_2S_2S_1_1440_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1314_in2 = bnn_Minus_2S_2S_1_1310_out1;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1314_in2 = bnn_Minus_2S_2S_1_1440_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_1308_ctrl1 or bnn_N_Mux_2_2_3_4_1314_in3 or bnn_N_Mux_2_2_3_4_1314_in2)
          begin :bnn_N_Mux_2_2_3_4_1314
            if (bnn_N_Mux_2_2_3_4_1308_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1314_out1 = bnn_N_Mux_2_2_3_4_1314_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1314_out1 = bnn_N_Mux_2_2_3_4_1314_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_1_1075_out1 or bnn_Add_4Sx2S_4S_1_1312_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1315_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1315_in2 = bnn_Add_4Sx2S_5S_1_1075_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1315_in2 = {bnn_Add_4Sx2S_4S_1_1312_out1[3], bnn_Add_4Sx2S_4S_1_1312_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1315_in2 = bnn_Add_4Sx2S_5S_1_1075_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1315
         assign bnn_Add_5Sx4S_6S_1_1315_out1 = {bnn_Add_5Sx4S_6S_1_1315_in2[4], bnn_Add_5Sx4S_6S_1_1315_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1311_out1[1]}}, bnn_N_Mux_2_2_3_1_1311_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_65_mi61 or s_reg_1112 or s_reg_931 or bnn_N_Mux_2_2_3_1_2089_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1316_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1316_in1 = bnn_N_Mux_2_2_3_1_2089_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1316_in1 = Bline_buffer_65_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1316_in1 = s_reg_931;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1316
         assign bnn_Minus_2S_2S_4_1316_out1 = -bnn_Minus_2S_2S_4_1316_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1317
         assign bnn_Minus_2S_2S_4_1317_out1 = -bnn_Minus_2S_2S_4_1316_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_73_mi61 or s_reg_1112 or s_reg_961 or bnn_N_Mux_64_2_2_1_1636_out1[50] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1318_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1318_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[50], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1318_in1 = Bline_buffer_73_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1318_in1 = s_reg_961;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1318
         assign bnn_Minus_2S_2S_4_1318_out1 = -bnn_Minus_2S_2S_4_1318_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1319
         assign bnn_Minus_2S_2S_4_1319_out1 = -bnn_Minus_2S_2S_4_1318_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1320
         assign bnn_Minus_2S_2S_4_1320_out1 = -bnn_Minus_2S_2S_4_1318_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_65_mi61 or s_reg_1112 or s_reg_931 or bnn_N_Mux_2_2_3_1_2089_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1321_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1321_in3 = bnn_N_Mux_2_2_3_1_2089_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1321_in3 = Bline_buffer_65_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1321_in3 = s_reg_931;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_Minus_2S_2S_4_1316_out1 or bnn_N_Mux_2_2_3_4_1321_in3)
          begin :bnn_N_Mux_2_2_3_4_1321
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_1321_out1 = bnn_Minus_2S_2S_4_1316_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1321_out1 = bnn_N_Mux_2_2_3_4_1321_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_Minus_2S_2S_4_1317_out1 or bnn_N_Mux_2_2_3_4_1321_in3)
          begin :bnn_N_Mux_2_2_3_4_1322
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_1322_out1 = bnn_Minus_2S_2S_4_1317_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1322_out1 = bnn_N_Mux_2_2_3_4_1321_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_66_mi61 or s_reg_1112 or s_reg_938 or bnn_N_Mux_2_2_3_1_2106_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1323_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1323_in1 = bnn_N_Mux_2_2_3_1_2106_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1323_in1 = Bline_buffer_66_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1323_in1 = s_reg_938;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1323
         assign bnn_Minus_2S_2S_4_1323_out1 = -bnn_Minus_2S_2S_4_1323_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1324
         assign bnn_Minus_2S_2S_1_1324_out1 = -bnn_Minus_2S_2S_4_1323_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1325
         assign bnn_Minus_2S_2S_1_1325_out1 = -bnn_Minus_2S_2S_4_1316_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_73_mi61 or s_reg_1112 or s_reg_961 or bnn_N_Mux_64_2_2_1_1636_out1[50] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1326_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1326_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[50], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1326_in3 = Bline_buffer_73_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1326_in3 = s_reg_961;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1318_out1 or bnn_N_Mux_2_2_3_4_1326_in3)
          begin :bnn_N_Mux_2_2_3_4_1326
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1326_out1 = bnn_Minus_2S_2S_4_1318_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1326_out1 = bnn_N_Mux_2_2_3_4_1326_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_74_mi61 or s_reg_1112 or s_reg_964 or bnn_N_Mux_64_2_2_1_1636_out1[51] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1327_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1327_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[51], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1327_in1 = Bline_buffer_74_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1327_in1 = s_reg_964;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1327
         assign bnn_Minus_2S_2S_4_1327_out1 = -bnn_Minus_2S_2S_4_1327_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1319_out1 or bnn_N_Mux_2_2_3_4_1326_in3)
          begin :bnn_N_Mux_2_2_3_4_1328
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1328_out1 = bnn_Minus_2S_2S_4_1319_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1328_out1 = bnn_N_Mux_2_2_3_4_1326_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1329
         assign bnn_Minus_2S_2S_4_1329_out1 = -bnn_Minus_2S_2S_4_1327_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1320_out1 or bnn_N_Mux_2_2_3_4_1326_in3)
          begin :bnn_N_Mux_2_2_3_4_1330
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1330_out1 = bnn_Minus_2S_2S_4_1320_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1330_out1 = bnn_N_Mux_2_2_3_4_1326_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1331
         assign bnn_Add_3Sx3S_4S_4_1331_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1321_out1[1]}}, bnn_N_Mux_2_2_3_4_1321_out1} + {bnn_Add_2Sx2S_3S_4_1274_out1[2], bnn_Add_2Sx2S_3S_4_1274_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1332
         assign bnn_Minus_2S_2S_4_1332_out1 = -bnn_Minus_2S_2S_4_1327_in1;

         // resource: bnn_Add_2Sx2S_3S_4  instance: bnn_Add_2Sx2S_3S_4_1333
         assign bnn_Add_2Sx2S_3S_4_1333_out1 = {bnn_N_Mux_2_2_3_4_1279_out1[1], bnn_N_Mux_2_2_3_4_1279_out1} + {bnn_N_Mux_2_2_3_4_1322_out1[1], bnn_N_Mux_2_2_3_4_1322_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_66_mi61 or s_reg_1112 or s_reg_938 or bnn_N_Mux_2_2_3_1_2106_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1334_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1334_in3 = bnn_N_Mux_2_2_3_1_2106_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1334_in3 = Bline_buffer_66_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1334_in3 = s_reg_938;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_Minus_2S_2S_4_1323_out1 or bnn_N_Mux_2_2_3_4_1334_in3)
          begin :bnn_N_Mux_2_2_3_4_1334
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_1334_out1 = bnn_Minus_2S_2S_4_1323_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1334_out1 = bnn_N_Mux_2_2_3_4_1334_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_Minus_2S_2S_1_1324_out1 or bnn_N_Mux_2_2_3_4_1334_in3)
          begin :bnn_N_Mux_2_2_3_1_1335
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1335_out1 = bnn_Minus_2S_2S_1_1324_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1335_out1 = bnn_N_Mux_2_2_3_4_1334_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_4_1321_in3 or bnn_Minus_2S_2S_1_1325_out1)
          begin :bnn_N_Mux_2_2_3_1_1336
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1336_out1 = bnn_Minus_2S_2S_1_1325_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1336_out1 = bnn_N_Mux_2_2_3_4_1321_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1337
         assign bnn_Minus_2S_2S_1_1337_out1 = -bnn_Minus_2S_2S_4_1284_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1338
         assign bnn_Minus_2S_2S_1_1338_out1 = -bnn_Minus_2S_2S_4_1284_in1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1339
         assign bnn_Minus_2S_2S_1_1339_out1 = -bnn_Minus_2S_2S_4_1323_in1;

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_1340
         assign bnn_Add_4Sx2S_5S_1_1340_out1 = {bnn_Add_4Sx2S_4S_1_1281_out1[3], bnn_Add_4Sx2S_4S_1_1281_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1326_out1[1]}}, bnn_N_Mux_2_2_3_4_1326_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_74_mi61 or s_reg_1112 or s_reg_964 or bnn_N_Mux_64_2_2_1_1636_out1[51] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1341_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1341_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[51], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1341_in3 = Bline_buffer_74_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1341_in3 = s_reg_964;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1327_out1 or bnn_N_Mux_2_2_3_4_1341_in3)
          begin :bnn_N_Mux_2_2_3_4_1341
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1341_out1 = bnn_Minus_2S_2S_4_1327_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1341_out1 = bnn_N_Mux_2_2_3_4_1341_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1342
         assign bnn_Add_4Sx3S_4S_1_1342_out1 = bnn_Add_4Sx3S_4S_1_1282_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1328_out1[1]}}, bnn_N_Mux_2_2_3_4_1328_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_75_mi61 or s_reg_1112 or s_reg_967 or bnn_N_Mux_64_2_2_1_1636_out1[52] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1343_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1343_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[52], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1343_in1 = Bline_buffer_75_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1343_in1 = s_reg_967;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1343
         assign bnn_Minus_2S_2S_4_1343_out1 = -bnn_Minus_2S_2S_4_1343_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1329_out1 or bnn_N_Mux_2_2_3_4_1341_in3)
          begin :bnn_N_Mux_2_2_3_4_1344
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1344_out1 = bnn_Minus_2S_2S_4_1329_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1344_out1 = bnn_N_Mux_2_2_3_4_1341_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1345
         assign bnn_Add_4Sx2S_5S_4_1345_out1 = {bnn_Add_3Sx3S_4S_4_1331_out1[3], bnn_Add_3Sx3S_4S_4_1331_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1330_out1[1]}}, bnn_N_Mux_2_2_3_4_1330_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1346
         assign bnn_Minus_2S_2S_4_1346_out1 = -bnn_Minus_2S_2S_4_1343_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_1332_out1 or bnn_N_Mux_2_2_3_4_1341_in3)
          begin :bnn_N_Mux_2_2_3_4_1347
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_1347_out1 = bnn_Minus_2S_2S_4_1332_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1347_out1 = bnn_N_Mux_2_2_3_4_1341_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1348
         assign bnn_Add_3Sx3S_4S_4_1348_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1334_out1[1]}}, bnn_N_Mux_2_2_3_4_1334_out1} + {bnn_Add_2Sx2S_3S_4_1333_out1[2], bnn_Add_2Sx2S_3S_4_1333_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1349
         assign bnn_Minus_2S_2S_1_1349_out1 = -bnn_Minus_2S_2S_4_1343_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1350
         assign bnn_Add_2Sx2S_3S_1_1350_out1 = {bnn_N_Mux_2_2_3_1_1336_out1[1], bnn_N_Mux_2_2_3_1_1336_out1} + {bnn_N_Mux_2_2_3_1_1335_out1[1], bnn_N_Mux_2_2_3_1_1335_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_N_Mux_2_2_3_4_1286_in3 or bnn_Minus_2S_2S_1_1337_out1)
          begin :bnn_N_Mux_2_2_3_1_1351
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1351_out1 = bnn_Minus_2S_2S_1_1337_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1351_out1 = bnn_N_Mux_2_2_3_4_1286_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_4_1286_in3 or bnn_Minus_2S_2S_1_1338_out1)
          begin :bnn_N_Mux_2_2_3_1_1352
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1352_out1 = bnn_Minus_2S_2S_1_1338_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1352_out1 = bnn_N_Mux_2_2_3_4_1286_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_4_1334_in3 or bnn_Minus_2S_2S_1_1339_out1)
          begin :bnn_N_Mux_2_2_3_1_1353
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1353_out1 = bnn_Minus_2S_2S_1_1339_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1353_out1 = bnn_N_Mux_2_2_3_4_1334_in3;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1354
         assign bnn_Minus_2S_2S_1_1354_out1 = -bnn_Minus_2S_2S_4_1283_in1;

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1355
         assign bnn_Add_4Sx2S_5S_4_1355_out1 = {bnn_Add_4Sx3S_4S_1_1342_out1[3], bnn_Add_4Sx3S_4S_1_1342_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1341_out1[1]}}, bnn_N_Mux_2_2_3_4_1341_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_75_mi61 or s_reg_1112 or s_reg_967 or bnn_N_Mux_64_2_2_1_1636_out1[52] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1356_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1356_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[52], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1356_in3 = Bline_buffer_75_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1356_in3 = s_reg_967;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1343_out1 or bnn_N_Mux_2_2_3_4_1356_in3)
          begin :bnn_N_Mux_2_2_3_4_1356
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1356_out1 = bnn_Minus_2S_2S_4_1343_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1356_out1 = bnn_N_Mux_2_2_3_4_1356_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1357
         assign bnn_Add_4Sx2S_5S_4_1357_out1 = {bnn_Add_4Sx2S_5S_4_1345_out1[3], bnn_Add_4Sx2S_5S_4_1345_out1[3:0]} + {{ 3 {bnn_N_Mux_2_2_3_4_1344_out1[1]}}, bnn_N_Mux_2_2_3_4_1344_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_76_mi61 or s_reg_1112 or s_reg_970 or bnn_N_Mux_64_2_2_1_1636_out1[53] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1358_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1358_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[53], 1'b1};
               end
               else begin
                  bnn_Minus_2S_2S_4_1358_in1 = Bline_buffer_76_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1358_in1 = s_reg_970;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1358
         assign bnn_Minus_2S_2S_4_1358_out1 = -bnn_Minus_2S_2S_4_1358_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_1346_out1 or bnn_N_Mux_2_2_3_4_1356_in3)
          begin :bnn_N_Mux_2_2_3_4_1359
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_1359_out1 = bnn_Minus_2S_2S_4_1346_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1359_out1 = bnn_N_Mux_2_2_3_4_1356_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1360
         assign bnn_Add_4Sx2S_5S_4_1360_out1 = {bnn_Add_3Sx3S_4S_4_1348_out1[3], bnn_Add_3Sx3S_4S_4_1348_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_1347_out1[1]}}, bnn_N_Mux_2_2_3_4_1347_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1361
         assign bnn_Minus_2S_2S_1_1361_out1 = -bnn_Minus_2S_2S_4_1358_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1349_out1 or bnn_N_Mux_2_2_3_4_1356_in3)
          begin :bnn_N_Mux_2_2_3_1_1362
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1362_out1 = bnn_Minus_2S_2S_1_1349_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1362_out1 = bnn_N_Mux_2_2_3_4_1356_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1363
         assign bnn_Add_3Sx3S_4S_1_1363_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1351_out1[1]}}, bnn_N_Mux_2_2_3_1_1351_out1} + {bnn_Add_2Sx2S_3S_1_1350_out1[2], bnn_Add_2Sx2S_3S_1_1350_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1364
         assign bnn_Minus_2S_2S_1_1364_out1 = -bnn_Minus_2S_2S_4_1358_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1365
         assign bnn_Add_2Sx2S_3S_1_1365_out1 = {bnn_N_Mux_2_2_3_1_1353_out1[1], bnn_N_Mux_2_2_3_1_1353_out1} + {bnn_N_Mux_2_2_3_1_1352_out1[1], bnn_N_Mux_2_2_3_1_1352_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_N_Mux_2_2_3_4_1285_in3 or bnn_Minus_2S_2S_1_1354_out1)
          begin :bnn_N_Mux_2_2_3_1_1366
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_1366_out1 = bnn_Minus_2S_2S_1_1354_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1366_out1 = bnn_N_Mux_2_2_3_4_1285_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1367
         assign bnn_Add_4Sx2S_5S_4_1367_out1 = {bnn_Add_4Sx2S_5S_4_1357_out1[3], bnn_Add_4Sx2S_5S_4_1357_out1[3:0]} + {{ 3 {bnn_N_Mux_2_2_3_4_1356_out1[1]}}, bnn_N_Mux_2_2_3_4_1356_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_76_mi61 or s_reg_1112 or s_reg_970 or bnn_N_Mux_64_2_2_1_1636_out1[53] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1368_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1368_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[53], 1'b1};
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1368_in3 = Bline_buffer_76_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1368_in3 = s_reg_970;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_1358_out1 or bnn_N_Mux_2_2_3_4_1368_in3)
          begin :bnn_N_Mux_2_2_3_4_1368
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_1368_out1 = bnn_Minus_2S_2S_4_1358_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1368_out1 = bnn_N_Mux_2_2_3_4_1368_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1369
         assign bnn_Add_4Sx2S_5S_4_1369_out1 = {bnn_Add_4Sx2S_5S_4_1360_out1[3], bnn_Add_4Sx2S_5S_4_1360_out1[3:0]} + {{ 3 {bnn_N_Mux_2_2_3_4_1359_out1[1]}}, bnn_N_Mux_2_2_3_4_1359_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_1361_out1 or bnn_N_Mux_2_2_3_4_1368_in3)
          begin :bnn_N_Mux_2_2_3_1_1371
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_1371_out1 = bnn_Minus_2S_2S_1_1361_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1371_out1 = bnn_N_Mux_2_2_3_4_1368_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1372
         assign bnn_Add_4Sx2S_4S_1_1372_out1 = bnn_Add_3Sx3S_4S_1_1363_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1362_out1[1]}}, bnn_N_Mux_2_2_3_1_1362_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1373
         assign bnn_Minus_2S_2S_1_1373_out1 = -bnn_Minus_2S_2S_1_1290_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_1364_out1 or bnn_N_Mux_2_2_3_4_1368_in3)
          begin :bnn_N_Mux_2_2_3_1_1374
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_1374_out1 = bnn_Minus_2S_2S_1_1364_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1374_out1 = bnn_N_Mux_2_2_3_4_1368_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1375
         assign bnn_Add_3Sx3S_4S_1_1375_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1366_out1[1]}}, bnn_N_Mux_2_2_3_1_1366_out1} + {bnn_Add_2Sx2S_3S_1_1365_out1[2], bnn_Add_2Sx2S_3S_1_1365_out1};

         // resource: bnn_Add_4Sx2S_5S_4  instance: bnn_Add_4Sx2S_5S_4_1378
         assign bnn_Add_4Sx2S_5S_4_1378_out1 = {bnn_Add_4Sx2S_5S_4_1369_out1[3], bnn_Add_4Sx2S_5S_4_1369_out1[3:0]} + {{ 3 {bnn_N_Mux_2_2_3_4_1368_out1[1]}}, bnn_N_Mux_2_2_3_4_1368_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_77_mi61 or s_reg_1112 or s_reg_873 or s_reg_994 or bnn_N_Mux_2_2_3_1_3093_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1379_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1379_in3 = bnn_N_Mux_2_2_3_1_3093_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1379_in3 = Bline_buffer_77_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1379_in3 = s_reg_994;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1379_in3 = s_reg_873;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1290_out1 or bnn_N_Mux_2_2_3_4_1308_ctrl1 or bnn_N_Mux_2_2_3_1_1379_in3)
          begin :bnn_N_Mux_2_2_3_1_1379
            if (bnn_N_Mux_2_2_3_4_1308_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1379_out1 = bnn_Minus_2S_2S_1_1290_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1379_out1 = bnn_N_Mux_2_2_3_1_1379_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_1_1037_out1 or bnn_Add_4Sx2S_4S_1_1372_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1380_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1380_in2 = bnn_Add_4Sx2S_5S_1_1037_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1380_in2 = {bnn_Add_4Sx2S_4S_1_1372_out1[3], bnn_Add_4Sx2S_4S_1_1372_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1380_in2 = bnn_Add_4Sx2S_5S_1_1037_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_1_1371_out1 or bnn_N_Mux_2_2_3_1_3630_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1380_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1380_in1_slice = bnn_N_Mux_2_2_3_1_3630_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1380_in1_slice = bnn_N_Mux_2_2_3_1_1371_out1;
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1380_in1_slice = bnn_N_Mux_2_2_3_1_3630_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1380
         assign bnn_Add_5Sx4S_6S_1_1380_out1 = {bnn_Add_5Sx4S_6S_1_1380_in2[4], bnn_Add_5Sx4S_6S_1_1380_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_1380_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_1380_in1_slice};

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_932 or s_reg_944 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1382_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1382_ctrl1 = s_reg_944;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1382_ctrl1 = s_reg_932;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1382_ctrl1 = s_reg_944;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1373_out1 or bnn_N_Mux_2_2_3_1_1379_in3 or bnn_N_Mux_2_2_3_1_1382_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1382
            if (bnn_N_Mux_2_2_3_1_1382_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1382_out1 = bnn_Minus_2S_2S_1_1373_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1382_out1 = bnn_N_Mux_2_2_3_1_1379_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1383
         assign bnn_Add_4Sx2S_4S_1_1383_out1 = bnn_Add_3Sx3S_4S_1_1375_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1374_out1[1]}}, bnn_N_Mux_2_2_3_1_1374_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1293_ctrl1 or bnn_Minus_2S_2S_1_1295_out1 or bnn_N_Mux_2_2_3_1_1301_in3)
          begin :bnn_N_Mux_2_2_3_1_1384
            if (bnn_N_Mux_2_2_3_1_1293_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1384_out1 = bnn_Minus_2S_2S_1_1295_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1384_out1 = bnn_N_Mux_2_2_3_1_1301_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_91_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1288_out1)
          begin :bnn_N_Mux_2_2_3_1_1385
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1385_out1 = bnn_Minus_2S_2S_1_1288_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1385_out1 = Bline_buffer_91_mi61;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_93_mi61 or s_reg_1112 or s_reg_873 or s_reg_965 or bnn_N_Mux_2_2_3_1_3093_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1386_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1386_in1 = bnn_N_Mux_2_2_3_1_3093_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1386_in1 = Bline_buffer_93_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1386_in1 = s_reg_965;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1386_in1 = s_reg_873;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1386
         assign bnn_Minus_2S_2S_1_1386_out1 = -bnn_Minus_2S_2S_1_1386_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1380_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1389_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1389_in2 = bnn_Add_5Sx4S_6S_1_1380_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1389_in2 = {bnn_Add_5Sx4S_6S_1_1380_out1[3], bnn_Add_5Sx4S_6S_1_1380_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1389_in2 = bnn_Add_5Sx4S_6S_1_1380_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1389
         assign bnn_Add_5Sx4S_6S_1_1389_out1 = {bnn_Add_5Sx4S_6S_1_1389_in2[4], bnn_Add_5Sx4S_6S_1_1389_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1379_out1[1]}}, bnn_N_Mux_2_2_3_1_1379_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_78_mi61 or s_reg_1112 or s_reg_878 or s_reg_996 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1390_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1390_in3 = bnn_N_Mux_2_2_3_1_3114_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1390_in3 = Bline_buffer_78_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1390_in3 = s_reg_996;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1390_in3 = s_reg_878;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1296_out1 or bnn_N_Mux_2_2_3_4_1308_ctrl1 or bnn_N_Mux_2_2_3_1_1390_in3)
          begin :bnn_N_Mux_2_2_3_1_1390
            if (bnn_N_Mux_2_2_3_4_1308_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1390_out1 = bnn_Minus_2S_2S_1_1296_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1390_out1 = bnn_N_Mux_2_2_3_1_1390_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_1_1057_out1 or bnn_Add_4Sx2S_4S_1_1383_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1391_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1391_in2 = bnn_Add_4Sx2S_5S_1_1057_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1391_in2 = {bnn_Add_4Sx2S_4S_1_1383_out1[3], bnn_Add_4Sx2S_4S_1_1383_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1391_in2 = bnn_Add_4Sx2S_5S_1_1057_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1391
         assign bnn_Add_5Sx4S_6S_1_1391_out1 = {bnn_Add_5Sx4S_6S_1_1391_in2[4], bnn_Add_5Sx4S_6S_1_1391_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1382_out1[1]}}, bnn_N_Mux_2_2_3_1_1382_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_101_mi61 or s_reg_1112 or s_reg_895 or s_reg_982 or bnn_N_Mux_2_2_3_1_3229_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1392_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1392_in1 = bnn_N_Mux_2_2_3_1_3229_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1392_in1 = Bline_buffer_101_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1392_in1 = s_reg_982;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1392_in1 = s_reg_895;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1392
         assign bnn_Minus_2S_2S_1_1392_out1 = -bnn_Minus_2S_2S_1_1392_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1393
         assign bnn_Add_2Sx2S_3S_1_1393_out1 = {bnn_N_Mux_2_2_3_1_1385_out1[1], bnn_N_Mux_2_2_3_1_1385_out1} + {bnn_N_Mux_2_2_3_1_1384_out1[1], bnn_N_Mux_2_2_3_1_1384_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_93_mi61 or s_reg_1112 or s_reg_873 or bnn_N_Mux_2_2_3_1_3093_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1394_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1394_in3 = bnn_N_Mux_2_2_3_1_3093_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1394_in3 = Bline_buffer_93_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1394_in3 = s_reg_873;
            end
         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_916 or s_reg_957 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1394_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1394_ctrl1 = s_reg_957;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1394_ctrl1 = s_reg_916;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1394_ctrl1 = s_reg_957;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1386_out1 or bnn_N_Mux_2_2_3_1_1394_in3 or bnn_N_Mux_2_2_3_1_1394_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1394
            if (bnn_N_Mux_2_2_3_1_1394_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1394_out1 = bnn_Minus_2S_2S_1_1386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1394_out1 = bnn_N_Mux_2_2_3_1_1394_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_93_mi61 or s_reg_907 or bnn_Minus_2S_2S_1_1386_out1)
          begin :bnn_N_Mux_2_2_3_1_1395
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1395_out1 = bnn_Minus_2S_2S_1_1386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1395_out1 = Bline_buffer_93_mi61;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_92_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1295_out1)
          begin :bnn_N_Mux_2_2_3_1_1396
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1396_out1 = bnn_Minus_2S_2S_1_1295_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1396_out1 = Bline_buffer_92_mi61;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_94_mi61 or s_reg_1112 or s_reg_900 or s_reg_968 or bnn_N_Mux_2_2_3_1_3168_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1397_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1397_in1 = bnn_N_Mux_2_2_3_1_3168_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1397_in1 = Bline_buffer_94_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1397_in1 = s_reg_968;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1397_in1 = s_reg_900;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1397
         assign bnn_Minus_2S_2S_1_1397_out1 = -bnn_Minus_2S_2S_1_1397_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1391_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1400_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1400_in2 = bnn_Add_5Sx4S_6S_1_1391_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1400_in2 = {bnn_Add_5Sx4S_6S_1_1391_out1[3], bnn_Add_5Sx4S_6S_1_1391_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1400_in2 = bnn_Add_5Sx4S_6S_1_1391_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1400
         assign bnn_Add_5Sx4S_6S_1_1400_out1 = {bnn_Add_5Sx4S_6S_1_1400_in2[4], bnn_Add_5Sx4S_6S_1_1400_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1390_out1[1]}}, bnn_N_Mux_2_2_3_1_1390_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_101_mi61 or s_reg_1112 or s_reg_895 or s_reg_982 or bnn_N_Mux_2_2_3_1_3229_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1402_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1402_in3 = bnn_N_Mux_2_2_3_1_3229_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1402_in3 = Bline_buffer_101_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1402_in3 = s_reg_982;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1402_in3 = s_reg_895;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1392_out1 or bnn_N_Mux_2_2_3_1_1402_in3)
          begin :bnn_N_Mux_2_2_3_1_1402
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1402_out1 = bnn_Minus_2S_2S_1_1392_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1402_out1 = bnn_N_Mux_2_2_3_1_1402_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1403
         assign bnn_Add_3Sx3S_4S_1_1403_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1394_out1[1]}}, bnn_N_Mux_2_2_3_1_1394_out1} + {bnn_Add_2Sx2S_3S_1_1393_out1[2], bnn_Add_2Sx2S_3S_1_1393_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_102_mi61 or s_reg_1112 or s_reg_949 or bnn_N_Mux_2_2_3_1_3338_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_1_1404_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1404_in1 = bnn_N_Mux_2_2_3_1_3338_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1404_in1 = Bline_buffer_102_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1404_in1 = s_reg_949;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1404
         assign bnn_Minus_2S_2S_1_1404_out1 = -bnn_Minus_2S_2S_1_1404_in1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1405
         assign bnn_Add_2Sx2S_3S_1_1405_out1 = {bnn_N_Mux_2_2_3_1_1396_out1[1], bnn_N_Mux_2_2_3_1_1396_out1} + {bnn_N_Mux_2_2_3_1_1395_out1[1], bnn_N_Mux_2_2_3_1_1395_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_94_mi61 or s_reg_1112 or s_reg_900 or s_reg_968 or bnn_N_Mux_2_2_3_1_3168_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1406_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1406_in3 = bnn_N_Mux_2_2_3_1_3168_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1406_in3 = Bline_buffer_94_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1406_in3 = s_reg_968;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1406_in3 = s_reg_900;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_916 or s_reg_944 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1406_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1406_ctrl1 = s_reg_944;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1406_ctrl1 = s_reg_916;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1406_ctrl1 = s_reg_944;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1397_out1 or bnn_N_Mux_2_2_3_1_1406_in3 or bnn_N_Mux_2_2_3_1_1406_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1406
            if (bnn_N_Mux_2_2_3_1_1406_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1406_out1 = bnn_Minus_2S_2S_1_1397_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1406_out1 = bnn_N_Mux_2_2_3_1_1406_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_94_mi61 or s_reg_1112 or s_reg_900 or bnn_N_Mux_2_2_3_1_3168_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1407_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1407_in3 = bnn_N_Mux_2_2_3_1_3168_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1407_in3 = Bline_buffer_94_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1407_in3 = s_reg_900;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1293_ctrl1 or bnn_Minus_2S_2S_1_1397_out1 or bnn_N_Mux_2_2_3_1_1407_in3)
          begin :bnn_N_Mux_2_2_3_1_1407
            if (bnn_N_Mux_2_2_3_1_1293_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1407_out1 = bnn_Minus_2S_2S_1_1397_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1407_out1 = bnn_N_Mux_2_2_3_1_1407_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_93_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1386_out1)
          begin :bnn_N_Mux_2_2_3_1_1408
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1408_out1 = bnn_Minus_2S_2S_1_1386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1408_out1 = Bline_buffer_93_mi61;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_95_mi61 or s_reg_1112 or s_reg_878 or s_reg_971 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1409_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1409_in1 = bnn_N_Mux_2_2_3_1_3114_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1409_in1 = Bline_buffer_95_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1409_in1 = s_reg_971;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1409_in1 = s_reg_878;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1409
         assign bnn_Minus_2S_2S_1_1409_out1 = -bnn_Minus_2S_2S_1_1409_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_103_mi61 or s_reg_1112 or s_reg_904 or s_reg_986 or bnn_N_Mux_2_2_3_1_3243_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1418_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1418_in1 = bnn_N_Mux_2_2_3_1_3243_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1418_in1 = Bline_buffer_103_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1418_in1 = s_reg_986;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1418_in1 = s_reg_904;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1418
         assign bnn_Minus_2S_2S_1_1418_out1 = -bnn_Minus_2S_2S_1_1418_in1;

         // resource: mux_2bx4i
         always @(Bline_buffer_102_mi61 or s_reg_1112 or s_reg_895 or s_reg_982 or bnn_N_Mux_2_2_3_1_3229_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1413_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1413_in3 = bnn_N_Mux_2_2_3_1_3229_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1413_in3 = Bline_buffer_102_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1413_in3 = s_reg_982;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1413_in3 = s_reg_895;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_932 or s_reg_951 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1413_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1413_ctrl1 = s_reg_951;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1413_ctrl1 = s_reg_932;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1413_ctrl1 = s_reg_951;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1310_out1 or bnn_N_Mux_2_2_3_1_1413_in3 or bnn_N_Mux_2_2_3_1_1413_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1413
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1413_out1 = bnn_Minus_2S_2S_1_1310_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1413_out1 = bnn_N_Mux_2_2_3_1_1413_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1414
         assign bnn_Add_4Sx2S_4S_1_1414_out1 = bnn_Add_3Sx3S_4S_1_1403_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1402_out1[1]}}, bnn_N_Mux_2_2_3_1_1402_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_102_mi61 or s_reg_1112 or s_reg_949 or bnn_N_Mux_2_2_3_1_3338_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1416_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1416_in3 = bnn_N_Mux_2_2_3_1_3338_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1416_in3 = Bline_buffer_102_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1416_in3 = s_reg_949;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1404_out1 or bnn_N_Mux_2_2_3_1_1416_in3)
          begin :bnn_N_Mux_2_2_3_1_1416
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1416_out1 = bnn_Minus_2S_2S_1_1404_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1416_out1 = bnn_N_Mux_2_2_3_1_1416_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1417
         assign bnn_Add_3Sx3S_4S_1_1417_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1406_out1[1]}}, bnn_N_Mux_2_2_3_1_1406_out1} + {bnn_Add_2Sx2S_3S_1_1405_out1[2], bnn_Add_2Sx2S_3S_1_1405_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1419
         assign bnn_Add_2Sx2S_3S_1_1419_out1 = {bnn_N_Mux_2_2_3_1_1408_out1[1], bnn_N_Mux_2_2_3_1_1408_out1} + {bnn_N_Mux_2_2_3_1_1407_out1[1], bnn_N_Mux_2_2_3_1_1407_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_95_mi61 or s_reg_1112 or s_reg_878 or bnn_N_Mux_2_2_3_1_3114_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1420_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1420_in3 = bnn_N_Mux_2_2_3_1_3114_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1420_in3 = Bline_buffer_95_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1420_in3 = s_reg_878;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1394_ctrl1 or bnn_Minus_2S_2S_1_1409_out1 or bnn_N_Mux_2_2_3_1_1420_in3)
          begin :bnn_N_Mux_2_2_3_1_1420
            if (bnn_N_Mux_2_2_3_1_1394_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1420_out1 = bnn_Minus_2S_2S_1_1409_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1420_out1 = bnn_N_Mux_2_2_3_1_1420_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_95_mi61 or s_reg_907 or bnn_Minus_2S_2S_1_1409_out1)
          begin :bnn_N_Mux_2_2_3_1_1421
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1421_out1 = bnn_Minus_2S_2S_1_1409_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1421_out1 = Bline_buffer_95_mi61;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_94_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1397_out1)
          begin :bnn_N_Mux_2_2_3_1_1422
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1422_out1 = bnn_Minus_2S_2S_1_1397_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1422_out1 = Bline_buffer_94_mi61;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_96_mi61 or s_reg_1112 or s_reg_894 or s_reg_974 or bnn_N_Mux_2_2_3_1_3203_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1423_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1423_in1 = bnn_N_Mux_2_2_3_1_3203_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1423_in1 = Bline_buffer_96_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1423_in1 = s_reg_974;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1423_in1 = s_reg_894;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1423
         assign bnn_Minus_2S_2S_1_1423_out1 = -bnn_Minus_2S_2S_1_1423_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1315_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_4_1426_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_4_1426_in2 = bnn_Add_5Sx4S_6S_1_1315_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_4_1426_in2 = {bnn_Add_5Sx4S_6S_1_1315_out1[3], bnn_Add_5Sx4S_6S_1_1315_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_4_1426_in2 = bnn_Add_5Sx4S_6S_1_1315_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1426
         assign bnn_Add_5Sx4S_6S_4_1426_out1 = {bnn_Add_5Sx4S_6S_4_1426_in2[4], bnn_Add_5Sx4S_6S_4_1426_in2} + {{ 4 {bnn_N_Mux_2_2_3_4_1314_out1[1]}}, bnn_N_Mux_2_2_3_4_1314_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_103_mi61 or s_reg_1112 or s_reg_904 or s_reg_986 or bnn_N_Mux_2_2_3_1_3243_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1427_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1427_in3 = bnn_N_Mux_2_2_3_1_3243_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1427_in3 = Bline_buffer_103_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1427_in3 = s_reg_986;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1427_in3 = s_reg_904;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(s_reg_1112 or s_reg_939 or s_reg_957 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1427_ctrl1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1427_ctrl1 = s_reg_957;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1427_ctrl1 = s_reg_939;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1427_ctrl1 = s_reg_957;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1418_out1 or bnn_N_Mux_2_2_3_1_1427_in3 or bnn_N_Mux_2_2_3_1_1427_ctrl1)
          begin :bnn_N_Mux_2_2_3_1_1427
            if (bnn_N_Mux_2_2_3_1_1427_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1427_out1 = bnn_Minus_2S_2S_1_1418_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1427_out1 = bnn_N_Mux_2_2_3_1_1427_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_6Ux6U_6U_1_274_out1[4:0] or bnn_Add_4Sx2S_4S_1_1414_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1428_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1428_in2 = bnn_Add_6Ux6U_6U_1_274_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1428_in2 = {bnn_Add_4Sx2S_4S_1_1414_out1[3], bnn_Add_4Sx2S_4S_1_1414_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1428_in2 = bnn_Add_6Ux6U_6U_1_274_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1428
         assign bnn_Add_5Sx4S_6S_1_1428_out1 = {bnn_Add_5Sx4S_6S_1_1428_in2[4], bnn_Add_5Sx4S_6S_1_1428_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1413_out1[1]}}, bnn_N_Mux_2_2_3_1_1413_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_104_mi61 or s_reg_1112 or s_reg_914 or s_reg_988 or bnn_N_Mux_2_2_3_1_3258_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1435_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1435_in1 = bnn_N_Mux_2_2_3_1_3258_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1435_in1 = Bline_buffer_104_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1435_in1 = s_reg_988;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1435_in1 = s_reg_914;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1435
         assign bnn_Minus_2S_2S_1_1435_out1 = -bnn_Minus_2S_2S_1_1435_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Minus_2S_2S_1_1418_out1 or bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_N_Mux_2_2_3_1_1427_in3)
          begin :bnn_N_Mux_2_2_3_1_1430
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1430_out1 = bnn_Minus_2S_2S_1_1418_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1430_out1 = bnn_N_Mux_2_2_3_1_1427_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1431
         assign bnn_Add_4Sx2S_4S_1_1431_out1 = bnn_Add_3Sx3S_4S_1_1417_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1416_out1[1]}}, bnn_N_Mux_2_2_3_1_1416_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1418_out1 or bnn_N_Mux_2_2_3_1_1427_in3)
          begin :bnn_N_Mux_2_2_3_1_1433
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1433_out1 = bnn_Minus_2S_2S_1_1418_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1433_out1 = bnn_N_Mux_2_2_3_1_1427_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1434
         assign bnn_Add_3Sx3S_4S_1_1434_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1420_out1[1]}}, bnn_N_Mux_2_2_3_1_1420_out1} + {bnn_Add_2Sx2S_3S_1_1419_out1[2], bnn_Add_2Sx2S_3S_1_1419_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1436
         assign bnn_Add_2Sx2S_3S_1_1436_out1 = {bnn_N_Mux_2_2_3_1_1422_out1[1], bnn_N_Mux_2_2_3_1_1422_out1} + {bnn_N_Mux_2_2_3_1_1421_out1[1], bnn_N_Mux_2_2_3_1_1421_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_96_mi61 or s_reg_1112 or s_reg_894 or bnn_N_Mux_2_2_3_1_3203_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_1437_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_1_1437_in3 = bnn_N_Mux_2_2_3_1_3203_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_1_1437_in3 = Bline_buffer_96_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_1_1437_in3 = s_reg_894;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1406_ctrl1 or bnn_Minus_2S_2S_1_1423_out1 or bnn_N_Mux_2_2_3_1_1437_in3)
          begin :bnn_N_Mux_2_2_3_1_1437
            if (bnn_N_Mux_2_2_3_1_1406_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1437_out1 = bnn_Minus_2S_2S_1_1423_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1437_out1 = bnn_N_Mux_2_2_3_1_1437_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_96_mi61 or s_reg_907 or bnn_Minus_2S_2S_1_1423_out1)
          begin :bnn_N_Mux_2_2_3_1_1438
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_1438_out1 = bnn_Minus_2S_2S_1_1423_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1438_out1 = Bline_buffer_96_mi61;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(Bline_buffer_95_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1409_out1)
          begin :bnn_N_Mux_2_2_3_1_1439
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_1439_out1 = bnn_Minus_2S_2S_1_1409_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1439_out1 = Bline_buffer_95_mi61;
            end
         end

         // resource: mux_2bx4i
         always @(Bline_buffer_97_mi61 or s_reg_1112 or s_reg_884 or s_reg_962 or bnn_N_Mux_2_2_3_1_3133_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1440_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1440_in1 = bnn_N_Mux_2_2_3_1_3133_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1440_in1 = Bline_buffer_97_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1440_in1 = s_reg_962;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1440_in1 = s_reg_884;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1440
         assign bnn_Minus_2S_2S_1_1440_out1 = -bnn_Minus_2S_2S_1_1440_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1428_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1443_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1443_in2 = bnn_Add_5Sx4S_6S_1_1428_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1443_in2 = {bnn_Add_5Sx4S_6S_1_1428_out1[3], bnn_Add_5Sx4S_6S_1_1428_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1443_in2 = bnn_Add_5Sx4S_6S_1_1428_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1443
         assign bnn_Add_5Sx4S_6S_1_1443_out1 = {bnn_Add_5Sx4S_6S_1_1443_in2[4], bnn_Add_5Sx4S_6S_1_1443_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1427_out1[1]}}, bnn_N_Mux_2_2_3_1_1427_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_104_mi61 or s_reg_1112 or s_reg_914 or s_reg_988 or bnn_N_Mux_2_2_3_1_3258_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1444_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1444_in3 = bnn_N_Mux_2_2_3_1_3258_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1444_in3 = Bline_buffer_104_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1444_in3 = s_reg_988;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1444_in3 = s_reg_914;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1427_ctrl1 or bnn_Minus_2S_2S_1_1435_out1 or bnn_N_Mux_2_2_3_1_1444_in3)
          begin :bnn_N_Mux_2_2_3_1_1444
            if (bnn_N_Mux_2_2_3_1_1427_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1444_out1 = bnn_Minus_2S_2S_1_1435_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1444_out1 = bnn_N_Mux_2_2_3_1_1444_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_6Ux6U_6U_1_314_out1[4:0] or bnn_Add_4Sx2S_4S_1_1431_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1445_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1445_in2 = bnn_Add_6Ux6U_6U_1_314_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1445_in2 = {bnn_Add_4Sx2S_4S_1_1431_out1[3], bnn_Add_4Sx2S_4S_1_1431_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1445_in2 = bnn_Add_6Ux6U_6U_1_314_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1445
         assign bnn_Add_5Sx4S_6S_1_1445_out1 = {bnn_Add_5Sx4S_6S_1_1445_in2[4], bnn_Add_5Sx4S_6S_1_1445_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1430_out1[1]}}, bnn_N_Mux_2_2_3_1_1430_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_105_mi61 or s_reg_1112 or s_reg_922 or s_reg_990 or bnn_N_Mux_2_2_3_1_3274_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1452_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1452_in1 = bnn_N_Mux_2_2_3_1_3274_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1452_in1 = Bline_buffer_105_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1452_in1 = s_reg_990;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1452_in1 = s_reg_922;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1452
         assign bnn_Minus_2S_2S_1_1452_out1 = -bnn_Minus_2S_2S_1_1452_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_Minus_2S_2S_1_1435_out1 or bnn_N_Mux_2_2_3_1_1444_in3)
          begin :bnn_N_Mux_2_2_3_1_1447
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1447_out1 = bnn_Minus_2S_2S_1_1435_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1447_out1 = bnn_N_Mux_2_2_3_1_1444_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1448
         assign bnn_Add_4Sx2S_4S_1_1448_out1 = bnn_Add_3Sx3S_4S_1_1434_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1433_out1[1]}}, bnn_N_Mux_2_2_3_1_1433_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1435_out1 or bnn_N_Mux_2_2_3_1_1444_in3)
          begin :bnn_N_Mux_2_2_3_1_1450
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1450_out1 = bnn_Minus_2S_2S_1_1435_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1450_out1 = bnn_N_Mux_2_2_3_1_1444_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1451
         assign bnn_Add_3Sx3S_4S_1_1451_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1437_out1[1]}}, bnn_N_Mux_2_2_3_1_1437_out1} + {bnn_Add_2Sx2S_3S_1_1436_out1[2], bnn_Add_2Sx2S_3S_1_1436_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1453
         assign bnn_Add_2Sx2S_3S_1_1453_out1 = {bnn_N_Mux_2_2_3_1_1439_out1[1], bnn_N_Mux_2_2_3_1_1439_out1} + {bnn_N_Mux_2_2_3_1_1438_out1[1], bnn_N_Mux_2_2_3_1_1438_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_97_mi61 or s_reg_1112 or s_reg_884 or s_reg_962 or bnn_N_Mux_2_2_3_1_3133_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1454_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1454_in3 = bnn_N_Mux_2_2_3_1_3133_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1454_in3 = Bline_buffer_97_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1454_in3 = s_reg_962;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1454_in3 = s_reg_884;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1406_ctrl1 or bnn_Minus_2S_2S_1_1440_out1 or bnn_N_Mux_2_2_3_1_1454_in3)
          begin :bnn_N_Mux_2_2_3_1_1454
            if (bnn_N_Mux_2_2_3_1_1406_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1454_out1 = bnn_Minus_2S_2S_1_1440_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1454_out1 = bnn_N_Mux_2_2_3_1_1454_in3;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_97_mi61 or s_reg_1112 or s_reg_884 or bnn_N_Mux_2_2_3_1_3133_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1455_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1455_in3 = bnn_N_Mux_2_2_3_1_3133_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1455_in3 = Bline_buffer_97_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1455_in3 = s_reg_884;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1293_ctrl1 or bnn_Minus_2S_2S_1_1440_out1 or bnn_N_Mux_2_2_3_4_1455_in3)
          begin :bnn_N_Mux_2_2_3_4_1455
            if (bnn_N_Mux_2_2_3_1_1293_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1455_out1 = bnn_Minus_2S_2S_1_1440_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1455_out1 = bnn_N_Mux_2_2_3_4_1455_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(Bline_buffer_96_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1423_out1)
          begin :bnn_N_Mux_2_2_3_4_1456
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1456_out1 = bnn_Minus_2S_2S_1_1423_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1456_out1 = Bline_buffer_96_mi61;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_98_mi61 or s_reg_1112 or s_reg_919 or bnn_N_Mux_2_2_3_4_3200_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Minus_2S_2S_4_1457_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1457_in1 = bnn_N_Mux_2_2_3_4_3200_out1;
               end
               else begin
                  bnn_Minus_2S_2S_4_1457_in1 = Bline_buffer_98_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1457_in1 = s_reg_919;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1457
         assign bnn_Minus_2S_2S_4_1457_out1 = -bnn_Minus_2S_2S_4_1457_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1445_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1460_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1460_in2 = bnn_Add_5Sx4S_6S_1_1445_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1460_in2 = {bnn_Add_5Sx4S_6S_1_1445_out1[3], bnn_Add_5Sx4S_6S_1_1445_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1460_in2 = bnn_Add_5Sx4S_6S_1_1445_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1460
         assign bnn_Add_5Sx4S_6S_1_1460_out1 = {bnn_Add_5Sx4S_6S_1_1460_in2[4], bnn_Add_5Sx4S_6S_1_1460_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1444_out1[1]}}, bnn_N_Mux_2_2_3_1_1444_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_105_mi61 or s_reg_1112 or s_reg_922 or s_reg_990 or bnn_N_Mux_2_2_3_1_3274_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1461_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1461_in3 = bnn_N_Mux_2_2_3_1_3274_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1461_in3 = Bline_buffer_105_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1461_in3 = s_reg_990;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1461_in3 = s_reg_922;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1427_ctrl1 or bnn_Minus_2S_2S_1_1452_out1 or bnn_N_Mux_2_2_3_1_1461_in3)
          begin :bnn_N_Mux_2_2_3_1_1461
            if (bnn_N_Mux_2_2_3_1_1427_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1461_out1 = bnn_Minus_2S_2S_1_1452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1461_out1 = bnn_N_Mux_2_2_3_1_1461_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_6Ux6U_6U_1_407_out1[4:0] or bnn_Add_4Sx2S_4S_1_1448_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1462_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1462_in2 = bnn_Add_6Ux6U_6U_1_407_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1462_in2 = {bnn_Add_4Sx2S_4S_1_1448_out1[3], bnn_Add_4Sx2S_4S_1_1448_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1462_in2 = bnn_Add_6Ux6U_6U_1_407_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1462
         assign bnn_Add_5Sx4S_6S_1_1462_out1 = {bnn_Add_5Sx4S_6S_1_1462_in2[4], bnn_Add_5Sx4S_6S_1_1462_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1447_out1[1]}}, bnn_N_Mux_2_2_3_1_1447_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_106_mi61 or s_reg_1112 or s_reg_930 or s_reg_992 or bnn_N_Mux_2_2_3_1_3290_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1469_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1469_in1 = bnn_N_Mux_2_2_3_1_3290_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1469_in1 = Bline_buffer_106_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1469_in1 = s_reg_992;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1469_in1 = s_reg_930;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1469
         assign bnn_Minus_2S_2S_1_1469_out1 = -bnn_Minus_2S_2S_1_1469_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_Minus_2S_2S_1_1452_out1 or bnn_N_Mux_2_2_3_1_1461_in3)
          begin :bnn_N_Mux_2_2_3_1_1464
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1464_out1 = bnn_Minus_2S_2S_1_1452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1464_out1 = bnn_N_Mux_2_2_3_1_1461_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1465
         assign bnn_Add_4Sx2S_4S_1_1465_out1 = bnn_Add_3Sx3S_4S_1_1451_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1450_out1[1]}}, bnn_N_Mux_2_2_3_1_1450_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1452_out1 or bnn_N_Mux_2_2_3_1_1461_in3)
          begin :bnn_N_Mux_2_2_3_1_1467
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1467_out1 = bnn_Minus_2S_2S_1_1452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1467_out1 = bnn_N_Mux_2_2_3_1_1461_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_1468
         assign bnn_Add_3Sx3S_4S_1_1468_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_1454_out1[1]}}, bnn_N_Mux_2_2_3_1_1454_out1} + {bnn_Add_2Sx2S_3S_1_1453_out1[2], bnn_Add_2Sx2S_3S_1_1453_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_1470
         assign bnn_Add_2Sx2S_3S_1_1470_out1 = {bnn_N_Mux_2_2_3_4_1456_out1[1], bnn_N_Mux_2_2_3_4_1456_out1} + {bnn_N_Mux_2_2_3_4_1455_out1[1], bnn_N_Mux_2_2_3_4_1455_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_98_mi61 or s_reg_1112 or s_reg_919 or bnn_N_Mux_2_2_3_4_3200_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1471_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1471_in3 = bnn_N_Mux_2_2_3_4_3200_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1471_in3 = Bline_buffer_98_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1471_in3 = s_reg_919;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_1292_ctrl1 or bnn_Minus_2S_2S_4_1457_out1 or bnn_N_Mux_2_2_3_4_1471_in3)
          begin :bnn_N_Mux_2_2_3_4_1471
            if (bnn_N_Mux_2_2_3_4_1292_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1471_out1 = bnn_Minus_2S_2S_4_1457_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1471_out1 = bnn_N_Mux_2_2_3_4_1471_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1293_ctrl1 or bnn_Minus_2S_2S_4_1457_out1 or bnn_N_Mux_2_2_3_4_1471_in3)
          begin :bnn_N_Mux_2_2_3_4_1472
            if (bnn_N_Mux_2_2_3_1_1293_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1472_out1 = bnn_Minus_2S_2S_4_1457_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1472_out1 = bnn_N_Mux_2_2_3_4_1471_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(Bline_buffer_97_mi61 or s_reg_908 or bnn_Minus_2S_2S_1_1440_out1)
          begin :bnn_N_Mux_2_2_3_4_1473
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1473_out1 = bnn_Minus_2S_2S_1_1440_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1473_out1 = Bline_buffer_97_mi61;
            end
         end

         // resource: mux_2bx3i
         always @(Bline_buffer_99_mi61 or s_reg_1112 or s_reg_883 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_2178_out1_slice)
          begin :drive_bnn_Minus_2S_2S_4_1474_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_4_1474_in1 = bnn_N_Mux_3_2_6_4_2178_out1_slice;
               end
               else begin
                  bnn_Minus_2S_2S_4_1474_in1 = Bline_buffer_99_mi61;
               end
            end
            else begin
               bnn_Minus_2S_2S_4_1474_in1 = s_reg_883;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_1474
         assign bnn_Minus_2S_2S_4_1474_out1 = -bnn_Minus_2S_2S_4_1474_in1;

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1462_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1475_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1475_in2 = bnn_Add_5Sx4S_6S_1_1462_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1475_in2 = {bnn_Add_5Sx4S_6S_1_1462_out1[3], bnn_Add_5Sx4S_6S_1_1462_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1475_in2 = bnn_Add_5Sx4S_6S_1_1462_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1475
         assign bnn_Add_5Sx4S_6S_1_1475_out1 = {bnn_Add_5Sx4S_6S_1_1475_in2[4], bnn_Add_5Sx4S_6S_1_1475_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1461_out1[1]}}, bnn_N_Mux_2_2_3_1_1461_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_106_mi61 or s_reg_1112 or s_reg_930 or s_reg_992 or bnn_N_Mux_2_2_3_1_3290_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1476_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1476_in3 = bnn_N_Mux_2_2_3_1_3290_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1476_in3 = Bline_buffer_106_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1476_in3 = s_reg_992;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1476_in3 = s_reg_930;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1427_ctrl1 or bnn_Minus_2S_2S_1_1469_out1 or bnn_N_Mux_2_2_3_1_1476_in3)
          begin :bnn_N_Mux_2_2_3_1_1476
            if (bnn_N_Mux_2_2_3_1_1427_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1476_out1 = bnn_Minus_2S_2S_1_1469_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1476_out1 = bnn_N_Mux_2_2_3_1_1476_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_6Ux6U_6U_1_282_out1[4:0] or bnn_Add_4Sx2S_4S_1_1465_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1477_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1477_in2 = bnn_Add_6Ux6U_6U_1_282_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1477_in2 = {bnn_Add_4Sx2S_4S_1_1465_out1[3], bnn_Add_4Sx2S_4S_1_1465_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1477_in2 = bnn_Add_6Ux6U_6U_1_282_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1477
         assign bnn_Add_5Sx4S_6S_1_1477_out1 = {bnn_Add_5Sx4S_6S_1_1477_in2[4], bnn_Add_5Sx4S_6S_1_1477_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1464_out1[1]}}, bnn_N_Mux_2_2_3_1_1464_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_107_mi61 or s_reg_1112 or s_reg_937 or s_reg_994 or bnn_N_Mux_2_2_3_1_3306_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1478_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1478_in1 = bnn_N_Mux_2_2_3_1_3306_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1478_in1 = Bline_buffer_107_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1478_in1 = s_reg_994;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1478_in1 = s_reg_937;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1478
         assign bnn_Minus_2S_2S_1_1478_out1 = -bnn_Minus_2S_2S_1_1478_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_Minus_2S_2S_1_1469_out1 or bnn_N_Mux_2_2_3_1_1476_in3)
          begin :bnn_N_Mux_2_2_3_1_1479
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1479_out1 = bnn_Minus_2S_2S_1_1469_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1479_out1 = bnn_N_Mux_2_2_3_1_1476_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_1480
         assign bnn_Add_4Sx2S_4S_1_1480_out1 = bnn_Add_3Sx3S_4S_1_1468_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_1467_out1[1]}}, bnn_N_Mux_2_2_3_1_1467_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_106_mi61 or s_reg_1112 or s_reg_930 or bnn_N_Mux_2_2_3_1_3290_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1482_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1482_in3 = bnn_N_Mux_2_2_3_1_3290_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1482_in3 = Bline_buffer_106_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1482_in3 = s_reg_930;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1469_out1 or bnn_N_Mux_2_2_3_4_1482_in3)
          begin :bnn_N_Mux_2_2_3_4_1482
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1482_out1 = bnn_Minus_2S_2S_1_1469_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1482_out1 = bnn_N_Mux_2_2_3_4_1482_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1483
         assign bnn_Add_3Sx3S_4S_4_1483_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1471_out1[1]}}, bnn_N_Mux_2_2_3_4_1471_out1} + {bnn_Add_2Sx2S_3S_1_1470_out1[2], bnn_Add_2Sx2S_3S_1_1470_out1};

         // resource: bnn_Add_2Sx2S_3S_4  instance: bnn_Add_2Sx2S_3S_4_1485
         assign bnn_Add_2Sx2S_3S_4_1485_out1 = {bnn_N_Mux_2_2_3_4_1473_out1[1], bnn_N_Mux_2_2_3_4_1473_out1} + {bnn_N_Mux_2_2_3_4_1472_out1[1], bnn_N_Mux_2_2_3_4_1472_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_99_mi61 or s_reg_1112 or s_reg_883 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_2178_out1_slice)
          begin :drive_bnn_N_Mux_2_2_3_4_1486_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1486_in3 = bnn_N_Mux_3_2_6_4_2178_out1_slice;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1486_in3 = Bline_buffer_99_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1486_in3 = s_reg_883;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1406_ctrl1 or bnn_Minus_2S_2S_4_1474_out1 or bnn_N_Mux_2_2_3_4_1486_in3)
          begin :bnn_N_Mux_2_2_3_4_1486
            if (bnn_N_Mux_2_2_3_1_1406_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1486_out1 = bnn_Minus_2S_2S_4_1474_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1486_out1 = bnn_N_Mux_2_2_3_4_1486_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1477_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1487_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1487_in2 = bnn_Add_5Sx4S_6S_1_1477_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1487_in2 = {bnn_Add_5Sx4S_6S_1_1477_out1[3], bnn_Add_5Sx4S_6S_1_1477_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1487_in2 = bnn_Add_5Sx4S_6S_1_1477_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1487
         assign bnn_Add_5Sx4S_6S_1_1487_out1 = {bnn_Add_5Sx4S_6S_1_1487_in2[4], bnn_Add_5Sx4S_6S_1_1487_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1476_out1[1]}}, bnn_N_Mux_2_2_3_1_1476_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_107_mi61 or s_reg_1112 or s_reg_937 or s_reg_994 or bnn_N_Mux_2_2_3_1_3306_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_1488_in3
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_N_Mux_2_2_3_1_1488_in3 = bnn_N_Mux_2_2_3_1_3306_out1;
                  end
                  else begin
                     bnn_N_Mux_2_2_3_1_1488_in3 = Bline_buffer_107_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_1488_in3 = s_reg_994;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_1488_in3 = s_reg_937;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1427_ctrl1 or bnn_Minus_2S_2S_1_1478_out1 or bnn_N_Mux_2_2_3_1_1488_in3)
          begin :bnn_N_Mux_2_2_3_1_1488
            if (bnn_N_Mux_2_2_3_1_1427_ctrl1) begin
               bnn_N_Mux_2_2_3_1_1488_out1 = bnn_Minus_2S_2S_1_1478_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1488_out1 = bnn_N_Mux_2_2_3_1_1488_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_6Ux6U_6U_1_298_out1[4:0] or bnn_Add_4Sx2S_4S_1_1480_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1489_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1489_in2 = bnn_Add_6Ux6U_6U_1_298_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1489_in2 = {bnn_Add_4Sx2S_4S_1_1480_out1[3], bnn_Add_4Sx2S_4S_1_1480_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1489_in2 = bnn_Add_6Ux6U_6U_1_298_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1489
         assign bnn_Add_5Sx4S_6S_1_1489_out1 = {bnn_Add_5Sx4S_6S_1_1489_in2[4], bnn_Add_5Sx4S_6S_1_1489_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1479_out1[1]}}, bnn_N_Mux_2_2_3_1_1479_out1};

         // resource: mux_2bx4i
         always @(Bline_buffer_108_mi61 or s_reg_1112 or s_reg_890 or s_reg_965 or bnn_N_Mux_2_2_3_1_3151_out1 or cycle2_state or gs_ctrl196)
          begin :drive_bnn_Minus_2S_2S_1_1490_in1
            case (gs_ctrl196) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Minus_2S_2S_1_1490_in1 = bnn_N_Mux_2_2_3_1_3151_out1;
                  end
                  else begin
                     bnn_Minus_2S_2S_1_1490_in1 = Bline_buffer_108_mi61;
                  end
               end
               
               2'd2: begin
                  bnn_Minus_2S_2S_1_1490_in1 = s_reg_965;
               end
               
               default: begin
                  bnn_Minus_2S_2S_1_1490_in1 = s_reg_890;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1490
         assign bnn_Minus_2S_2S_1_1490_out1 = -bnn_Minus_2S_2S_1_1490_in1;

         // resource: mux_2bx3i
         always @(Bline_buffer_107_mi61 or s_reg_1112 or s_reg_937 or bnn_N_Mux_2_2_3_1_3306_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1491_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1491_in3 = bnn_N_Mux_2_2_3_1_3306_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1491_in3 = Bline_buffer_107_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1491_in3 = s_reg_937;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_Minus_2S_2S_1_1478_out1 or bnn_N_Mux_2_2_3_4_1491_in3)
          begin :bnn_N_Mux_2_2_3_4_1491
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1491_out1 = bnn_Minus_2S_2S_1_1478_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1491_out1 = bnn_N_Mux_2_2_3_4_1491_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_1492
         assign bnn_Add_4Sx3S_4S_1_1492_out1 = bnn_Add_3Sx3S_4S_4_1483_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_1482_out1[1]}}, bnn_N_Mux_2_2_3_4_1482_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1306_ctrl1 or bnn_Minus_2S_2S_1_1478_out1 or bnn_N_Mux_2_2_3_4_1491_in3)
          begin :bnn_N_Mux_2_2_3_4_1494
            if (bnn_N_Mux_2_2_3_1_1306_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1494_out1 = bnn_Minus_2S_2S_1_1478_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1494_out1 = bnn_N_Mux_2_2_3_4_1491_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_4  instance: bnn_Add_3Sx3S_4S_4_1495
         assign bnn_Add_3Sx3S_4S_4_1495_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_1486_out1[1]}}, bnn_N_Mux_2_2_3_4_1486_out1} + {bnn_Add_2Sx2S_3S_4_1485_out1[2], bnn_Add_2Sx2S_3S_4_1485_out1};

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1489_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1496_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1496_in2 = bnn_Add_5Sx4S_6S_1_1489_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1496_in2 = {bnn_Add_5Sx4S_6S_1_1489_out1[3], bnn_Add_5Sx4S_6S_1_1489_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1496_in2 = bnn_Add_5Sx4S_6S_1_1489_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1496
         assign bnn_Add_5Sx4S_6S_1_1496_out1 = {bnn_Add_5Sx4S_6S_1_1496_in2[4], bnn_Add_5Sx4S_6S_1_1496_in2} + {{ 4 {bnn_N_Mux_2_2_3_1_1488_out1[1]}}, bnn_N_Mux_2_2_3_1_1488_out1};

         // resource: mux_2bx3i
         always @(Bline_buffer_108_mi61 or s_reg_1112 or s_reg_890 or bnn_N_Mux_2_2_3_1_3151_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1497_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1497_in3 = bnn_N_Mux_2_2_3_1_3151_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1497_in3 = Bline_buffer_108_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1497_in3 = s_reg_890;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_1308_ctrl1 or bnn_Minus_2S_2S_1_1490_out1 or bnn_N_Mux_2_2_3_4_1497_in3)
          begin :bnn_N_Mux_2_2_3_4_1497
            if (bnn_N_Mux_2_2_3_4_1308_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1497_out1 = bnn_Minus_2S_2S_1_1490_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1497_out1 = bnn_N_Mux_2_2_3_4_1497_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_1_1092_out1 or bnn_Add_4Sx3S_4S_1_1492_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_4_1498_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_4_1498_in2 = bnn_Add_4Sx2S_5S_1_1092_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_4_1498_in2 = {bnn_Add_4Sx3S_4S_1_1492_out1[3], bnn_Add_4Sx3S_4S_1_1492_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_4_1498_in2 = bnn_Add_4Sx2S_5S_1_1092_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_1_1454_out1 or bnn_N_Mux_2_2_3_4_1491_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_4_1498_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_4_1498_in1_slice = bnn_N_Mux_2_2_3_1_1454_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_4_1498_in1_slice = bnn_N_Mux_2_2_3_4_1491_out1;
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_4_1498_in1_slice = bnn_N_Mux_2_2_3_1_1454_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1498
         assign bnn_Add_5Sx4S_6S_4_1498_out1 = {bnn_Add_5Sx4S_6S_4_1498_in2[4], bnn_Add_5Sx4S_6S_4_1498_in2} + {{ 4 {bnn_Add_5Sx4S_6S_4_1498_in1_slice[1]}}, bnn_Add_5Sx4S_6S_4_1498_in1_slice};

         // resource: mux_2bx3i
         always @(Bline_buffer_108_mi61 or s_reg_1112 or s_reg_900 or bnn_N_Mux_2_2_3_1_3168_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1499_in3
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1499_in3 = bnn_N_Mux_2_2_3_1_3168_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1499_in3 = Bline_buffer_108_mi61;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1499_in3 = s_reg_900;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_Minus_2S_2S_1_1397_out1 or bnn_Minus_2S_2S_1_1490_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_1499_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_N_Mux_2_2_3_4_1499_in2 = bnn_Minus_2S_2S_1_1397_out1;
               end
               else begin
                  bnn_N_Mux_2_2_3_4_1499_in2 = bnn_Minus_2S_2S_1_1490_out1;
               end
            end
            else begin
               bnn_N_Mux_2_2_3_4_1499_in2 = bnn_Minus_2S_2S_1_1397_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_1_1413_ctrl1 or bnn_N_Mux_2_2_3_4_1499_in3 or bnn_N_Mux_2_2_3_4_1499_in2)
          begin :bnn_N_Mux_2_2_3_4_1499
            if (bnn_N_Mux_2_2_3_1_1413_ctrl1) begin
               bnn_N_Mux_2_2_3_4_1499_out1 = bnn_N_Mux_2_2_3_4_1499_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1499_out1 = bnn_N_Mux_2_2_3_4_1499_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_4Sx2S_5S_4_1109_out1 or bnn_Add_3Sx3S_4S_4_1495_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1500_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1500_in2 = bnn_Add_4Sx2S_5S_4_1109_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1500_in2 = {bnn_Add_3Sx3S_4S_4_1495_out1[3], bnn_Add_3Sx3S_4S_4_1495_out1};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1500_in2 = bnn_Add_4Sx2S_5S_4_1109_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_4_1494_out1 or bnn_N_Mux_2_2_3_1_3730_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1500_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1500_in1_slice = bnn_N_Mux_2_2_3_1_3730_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1500_in1_slice = bnn_N_Mux_2_2_3_4_1494_out1;
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1500_in1_slice = bnn_N_Mux_2_2_3_1_3730_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1500
         assign bnn_Add_5Sx4S_6S_1_1500_out1 = {bnn_Add_5Sx4S_6S_1_1500_in2[4], bnn_Add_5Sx4S_6S_1_1500_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_1500_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_1500_in1_slice};

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_4_1498_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1501_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1501_in2 = bnn_Add_5Sx4S_6S_4_1498_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1501_in2 = {bnn_Add_5Sx4S_6S_4_1498_out1[3], bnn_Add_5Sx4S_6S_4_1498_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1501_in2 = bnn_Add_5Sx4S_6S_4_1498_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1501
         assign bnn_Add_5Sx4S_6S_1_1501_out1 = {bnn_Add_5Sx4S_6S_1_1501_in2[4], bnn_Add_5Sx4S_6S_1_1501_in2} + {{ 4 {bnn_N_Mux_2_2_3_4_1497_out1[1]}}, bnn_N_Mux_2_2_3_4_1497_out1};

         // resource: mux_5bx2i
         always @(s_reg_1112 or bnn_Add_5Sx4S_6S_1_1500_out1[4:0] or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1502_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1502_in2 = bnn_Add_5Sx4S_6S_1_1500_out1[4:0];
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1502_in2 = {bnn_Add_5Sx4S_6S_1_1500_out1[3], bnn_Add_5Sx4S_6S_1_1500_out1[3:0]};
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1502_in2 = bnn_Add_5Sx4S_6S_1_1500_out1[4:0];
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1502
         assign bnn_Add_5Sx4S_6S_1_1502_out1 = {bnn_Add_5Sx4S_6S_1_1502_in2[4], bnn_Add_5Sx4S_6S_1_1502_in2} + {{ 4 {bnn_N_Mux_2_2_3_4_1499_out1[1]}}, bnn_N_Mux_2_2_3_4_1499_out1};

         // resource: mux_2bx3i
         always @(s_reg_1112 or s_reg_943 or bnn_N_Mux_2_2_3_4_3325_out1 or cycle2_state or gs_ctrl197 or bnn_N_Mux_3_2_6_4_961_out1_slice)
          begin :drive_bnn_Minus_2S_2S_1_1503_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Minus_2S_2S_1_1503_in1 = bnn_N_Mux_2_2_3_4_3325_out1;
               end
               else begin
                  bnn_Minus_2S_2S_1_1503_in1 = bnn_N_Mux_3_2_6_4_961_out1_slice;
               end
            end
            else begin
               bnn_Minus_2S_2S_1_1503_in1 = s_reg_943;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_1503
         assign bnn_Minus_2S_2S_1_1503_out1 = -bnn_Minus_2S_2S_1_1503_in1;

         assign bnn_Or_1Sx1U_1S_4_1504_in1 = s_reg_871[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1504
         assign bnn_Or_1Sx1U_1S_4_1504_out1 = s_reg_1037 | bnn_Or_1Sx1U_1S_4_1504_in1;

         assign bnn_Or_1Sx1U_1S_4_1505_in1 = s_reg_1035[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1505
         assign bnn_Or_1Sx1U_1S_4_1505_out1 = s_reg_1038 | bnn_Or_1Sx1U_1S_4_1505_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_1506
         assign bnn_GreaterThan_6Sx4S_1U_4_1506_out1 = s_reg_1039[4] ^ s_reg_1039 > 5'd07;

         assign bnn_Or_1Sx1U_1S_4_1507_in1 = s_reg_1032[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1507
         assign bnn_Or_1Sx1U_1S_4_1507_out1 = s_reg_1040 | bnn_Or_1Sx1U_1S_4_1507_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_1508
         assign bnn_GreaterThan_6Sx4S_1U_4_1508_out1 = s_reg_1041[5] ^ s_reg_1041[5:0] > 6'd07;

         assign bnn_Or_1Sx1U_1S_4_1509_in1 = s_reg_1036[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1509
         assign bnn_Or_1Sx1U_1S_4_1509_out1 = s_reg_1042 | bnn_Or_1Sx1U_1S_4_1509_in1;

         assign bnn_Or_1Sx1U_1S_4_1510_in1 = s_reg_1021[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1510
         assign bnn_Or_1Sx1U_1S_4_1510_out1 = s_reg_1045 | bnn_Or_1Sx1U_1S_4_1510_in1;

         assign bnn_Or_1Sx1U_1S_4_1511_in1 = s_reg_1043[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1511
         assign bnn_Or_1Sx1U_1S_4_1511_out1 = s_reg_1049 | bnn_Or_1Sx1U_1S_4_1511_in1;

         assign bnn_Or_1Sx1U_1S_4_1512_in1 = s_reg_1046[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1512
         assign bnn_Or_1Sx1U_1S_4_1512_out1 = s_reg_1051 | bnn_Or_1Sx1U_1S_4_1512_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_1513
         assign bnn_GreaterThan_6Sx4S_1U_4_1513_out1 = s_reg_1027[4] ^ s_reg_1027 > 5'd07;

         assign bnn_Or_1Sx1U_1S_4_1514_in1 = s_reg_1047[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1514
         assign bnn_Or_1Sx1U_1S_4_1514_out1 = s_reg_1055 | bnn_Or_1Sx1U_1S_4_1514_in1;

         // resource: bnn_GreaterThan_6Sx4S_1U_4  instance: bnn_GreaterThan_6Sx4S_1U_4_1515
         assign bnn_GreaterThan_6Sx4S_1U_4_1515_out1 = s_reg_1058[5] ^ s_reg_1058[5:0] > 6'd07;

         assign bnn_Or_1Sx1U_1S_4_1516_in1 = s_reg_1031[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1516
         assign bnn_Or_1Sx1U_1S_4_1516_out1 = s_reg_1062 | bnn_Or_1Sx1U_1S_4_1516_in1;

         assign bnn_Or_1Sx1U_1S_4_1517_in1 = s_reg_1067[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1517
         assign bnn_Or_1Sx1U_1S_4_1517_out1 = s_reg_1069 | bnn_Or_1Sx1U_1S_4_1517_in1;

         assign bnn_Sub_8Sx2S_8S_4_1518_in2 = {s_reg_1076[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1518
         assign bnn_Sub_8Sx2S_8S_4_1518_out1 = bnn_Sub_8Sx2S_8S_4_1518_in2 - 8'd001;

         assign bnn_Or_1Sx1U_1S_4_1519_in1 = s_reg_1030[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1519
         assign bnn_Or_1Sx1U_1S_4_1519_out1 = s_reg_1065 | bnn_Or_1Sx1U_1S_4_1519_in1;

         assign bnn_Sub_8Sx2S_8S_4_1520_in2 = {s_reg_1036, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1520
         assign bnn_Sub_8Sx2S_8S_4_1520_out1 = bnn_Sub_8Sx2S_8S_4_1520_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1522_in2 = {s_reg_1029[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1522
         assign bnn_Sub_8Sx2S_8S_4_1522_out1 = bnn_Sub_8Sx2S_8S_4_1522_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1525_in2 = {s_reg_1030, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1525
         assign bnn_Sub_8Sx2S_8S_4_1525_out1 = bnn_Sub_8Sx2S_8S_4_1525_in2 - 8'd001;

         // resource: mux_6bx3i
         always @(s_reg_1036 or s_reg_1112 or bnn_Add_5Sx4S_6S_1_216_out1[4:0] or bnn_Mod_4Ux32U_7U_4_4577_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_1526_in2
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_6Ux6U_6U_1_1526_in2 = {bnn_Add_5Sx4S_6S_1_216_out1[4], bnn_Add_5Sx4S_6S_1_216_out1[4:0]};
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_1526_in2 = {s_reg_1036[4], s_reg_1036};
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_1526_in2 = bnn_Mod_4Ux32U_7U_4_4577_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_1526_in2 = {bnn_Add_5Sx4S_6S_1_216_out1[4], bnn_Add_5Sx4S_6S_1_216_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_4_4032_out1 or bnn_LeftShift_9Ux3U_7U_4_4576_out1[6:1] or cycle2_state or gs_ctrl242)
          begin :drive_bnn_Add_6Ux6U_6U_1_1526_in1
            case (gs_ctrl242) 

               2'd1: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     bnn_Add_6Ux6U_6U_1_1526_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_4032_out1[1]}}, bnn_N_Mux_2_2_3_4_4032_out1};
                  end
                  else begin
                     bnn_Add_6Ux6U_6U_1_1526_in1 = 6'd01;
                  end
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_1526_in1 = bnn_LeftShift_9Ux3U_7U_4_4576_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_1526_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_4032_out1[1]}}, bnn_N_Mux_2_2_3_4_4032_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_1526
         assign bnn_Add_6Ux6U_6U_1_1526_out1 = bnn_Add_6Ux6U_6U_1_1526_in2 + bnn_Add_6Ux6U_6U_1_1526_in1;

         assign bnn_Sub_8Sx2S_8S_4_1527_in2 = {s_reg_1021[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1527
         assign bnn_Sub_8Sx2S_8S_4_1527_out1 = bnn_Sub_8Sx2S_8S_4_1527_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1529_in2 = {s_reg_1093[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1529
         assign bnn_Sub_8Sx2S_8S_4_1529_out1 = bnn_Sub_8Sx2S_8S_4_1529_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1531_in2 = {s_reg_1043, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1531
         assign bnn_Sub_8Sx2S_8S_4_1531_out1 = bnn_Sub_8Sx2S_8S_4_1531_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1533_in2 = {s_reg_1031[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1533
         assign bnn_Sub_8Sx2S_8S_4_1533_out1 = bnn_Sub_8Sx2S_8S_4_1533_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1536_in2 = {s_reg_1039, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1536
         assign bnn_Sub_8Sx2S_8S_4_1536_out1 = bnn_Sub_8Sx2S_8S_4_1536_in2 - 8'd001;

         // resource: bnn_Sub_4Ux1U_4S_4  instance: bnn_Sub_4Ux1U_4S_4_1538
         assign bnn_Sub_4Ux1U_4S_4_1538_out1 = s_reg_1034[3:0] - 4'd01;

         assign bnn_Sub_8Sx2S_8S_4_1540_in2 = {s_reg_1027, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1540
         assign bnn_Sub_8Sx2S_8S_4_1540_out1 = bnn_Sub_8Sx2S_8S_4_1540_in2 - 8'd001;

         // resource: mux_5bx2i
         always @(s_reg_1039 or s_reg_1112 or bnn_Add_4Sx2S_5S_1_1340_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1542_in2
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1542_in2 = bnn_Add_4Sx2S_5S_1_1340_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1542_in2 = s_reg_1039;
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1542_in2 = bnn_Add_4Sx2S_5S_1_1340_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1112 or bnn_N_Mux_2_2_3_1_1416_out1 or cycle2_state or gs_ctrl197)
          begin :drive_bnn_Add_5Sx4S_6S_1_1542_in1
            if (gs_ctrl197) begin
               if (!cycle2_state && !s_reg_1112) begin
                  bnn_Add_5Sx4S_6S_1_1542_in1_slice = bnn_N_Mux_2_2_3_1_1416_out1;
               end
               else begin
                  bnn_Add_5Sx4S_6S_1_1542_in1_slice = 2'd1;
               end
            end
            else begin
               bnn_Add_5Sx4S_6S_1_1542_in1_slice = bnn_N_Mux_2_2_3_1_1416_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_1542
         assign bnn_Add_5Sx4S_6S_1_1542_out1 = {bnn_Add_5Sx4S_6S_1_1542_in2[4], bnn_Add_5Sx4S_6S_1_1542_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_1542_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_1542_in1_slice};

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1552
         assign bnn_Add_5Sx4S_6S_4_1552_out1 = {s_reg_1027[4], s_reg_1027} + 6'd01;

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1556
         assign bnn_Add_5Sx4S_6S_4_1556_out1 = {s_reg_1041[4], s_reg_1041[4:0]} + 6'd01;

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_1565
         assign bnn_Add_5Sx4S_6S_4_1565_out1 = {s_reg_1058[4], s_reg_1058[4:0]} + 6'd01;

         // resource: bnn_LessThan_10Ux32U_1U_4  instance: bnn_LessThan_10Ux32U_1U_4_1576
         assign bnn_LessThan_10Ux32U_1U_4_1576_out1 = {22'b0000000000000000000000, s_reg_1020} < s_reg_1000;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1577
         assign bnn_And_1Sx1U_1U_4_1577_out1 = s_reg_1044_stage1 & s_reg_1037_stage1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1578
         assign bnn_And_1Sx1U_1U_4_1578_out1 = s_reg_870_stage1 & s_reg_1038_stage1;

         assign bnn_Or_1Sx1U_1S_4_1579_in1 = s_reg_1039_stage1[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1579
         assign bnn_Or_1Sx1U_1S_4_1579_out1 = s_reg_1040_stage1 | bnn_Or_1Sx1U_1S_4_1579_in1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1580
         assign bnn_And_1Sx1U_1U_4_1580_out1 = s_reg_1048_stage1 & s_reg_1042_stage1;

         assign bnn_Or_1Sx1U_1S_4_1581_in1 = s_reg_1041_stage1_slice[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1581
         assign bnn_Or_1Sx1U_1S_4_1581_out1 = s_reg_1045_stage1 | bnn_Or_1Sx1U_1S_4_1581_in1;

         // resource: bnn_OrReduction_10U_1U_4  instance: bnn_OrReduction_10U_1U_4_1582
         assign bnn_OrReduction_10U_1U_4_1582_out1 = |s_reg_1034_stage1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1584
         assign bnn_And_1Sx1U_1U_4_1584_out1 = s_reg_1061_stage1 & s_reg_1055_stage1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1585
         assign bnn_And_1Sx1U_1U_4_1585_out1 = s_reg_1063_stage1 & s_reg_1062_stage1;

         assign bnn_Or_1Sx1U_1S_4_1586_in1 = s_reg_1027_stage1[4];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1586
         assign bnn_Or_1Sx1U_1S_4_1586_out1 = s_reg_1064_stage1 | bnn_Or_1Sx1U_1S_4_1586_in1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1587
         assign bnn_And_1Sx1U_1U_4_1587_out1 = s_reg_1066_stage1 & s_reg_1065_stage1;

         assign bnn_Or_1Sx1U_1S_4_1588_in1 = s_reg_1058_stage1_slice[5];

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_1588
         assign bnn_Or_1Sx1U_1S_4_1588_out1 = s_reg_1012[0] | bnn_Or_1Sx1U_1S_4_1588_in1;

         assign bnn_Sub_8Sx2S_8S_4_1596_in2 = {s_reg_1046_stage1_slice, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1596
         assign bnn_Sub_8Sx2S_8S_4_1596_out1 = bnn_Sub_8Sx2S_8S_4_1596_in2 - 8'd001;

         // resource: bnn_Sub_4Ux1U_4S_4  instance: bnn_Sub_4Ux1U_4S_4_1597
         assign bnn_Sub_4Ux1U_4S_4_1597_out1 = s_reg_1034_stage1[3:0] - 4'd01;

         assign bnn_Sub_8Sx2S_8S_4_1600_in2 = {s_reg_1041_stage1_slice[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1600
         assign bnn_Sub_8Sx2S_8S_4_1600_out1 = bnn_Sub_8Sx2S_8S_4_1600_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1606_in2 = {s_reg_1047_stage1, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1606
         assign bnn_Sub_8Sx2S_8S_4_1606_out1 = bnn_Sub_8Sx2S_8S_4_1606_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1610_in2 = {s_reg_1058_stage1_slice[4:0], 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1610
         assign bnn_Sub_8Sx2S_8S_4_1610_out1 = bnn_Sub_8Sx2S_8S_4_1610_in2 - 8'd001;

         assign bnn_Sub_8Sx2S_8S_4_1619_in2 = {s_reg_1067_stage1_slice, 3'd0};

         // resource: bnn_Sub_8Sx2S_8S_4  instance: bnn_Sub_8Sx2S_8S_4_1619
         assign bnn_Sub_8Sx2S_8S_4_1619_out1 = bnn_Sub_8Sx2S_8S_4_1619_in2 - 8'd001;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_1630
         assign bnn_And_1Sx1U_1U_4_1630_out1 = s_reg_1111_stage1 & s_reg_1082;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_883 or s_reg_887 or s_reg_908)
          begin :bnn_N_Mux_2_2_3_4_1634
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_1634_out1 = s_reg_887;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1634_out1 = s_reg_883;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1033 or s_reg_957 or s_reg_977)
          begin :bnn_N_Mux_2_2_3_4_1635
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_1635_out1 = s_reg_1033;
            end
            else begin
               bnn_N_Mux_2_2_3_4_1635_out1 = s_reg_977;
            end
         end

         // resource: bnn_N_Mux_64_2_2_1
         always @(memresp_data[63:0] or memresp_m_stall_reg_full or memresp_m_stall_reg_slice)
          begin :bnn_N_Mux_64_2_2_1_1636
            if (memresp_m_stall_reg_full) begin
               bnn_N_Mux_64_2_2_1_1636_out1 = memresp_m_stall_reg_slice;
            end
            else begin
               bnn_N_Mux_64_2_2_1_1636_out1 = memresp_data[63:0];
            end
         end

         assign bnn_N_Mux_3_2_6_4_1637_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[40], bnn_N_Mux_64_2_2_1_1636_out1[40]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_1637_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_1637
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_1637_out1_slice = bnn_N_Mux_3_2_6_4_1637_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_1637_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_4_1638_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[39], bnn_N_Mux_64_2_2_1_1636_out1[39]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_1638_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_1638
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_1638_out1_slice = bnn_N_Mux_3_2_6_4_1638_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_1638_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_1_1639_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[48], bnn_N_Mux_64_2_2_1_1636_out1[48]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1639_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1639
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1639_out1_slice = bnn_N_Mux_3_2_6_1_1639_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1639_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_4_1640_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[47], bnn_N_Mux_64_2_2_1_1636_out1[47]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_N_Mux_3_2_6_4_1640_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_4_1640
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_4_1640_out1_slice = bnn_N_Mux_3_2_6_4_1640_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_1640_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_1_1641_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[56], bnn_N_Mux_64_2_2_1_1636_out1[56]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1641_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1641
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1641_out1_slice = bnn_N_Mux_3_2_6_1_1641_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1641_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_1_1642_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[55], bnn_N_Mux_64_2_2_1_1636_out1[55]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1642_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1642
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1642_out1_slice = bnn_N_Mux_3_2_6_1_1642_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1642_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1643_in1 = {s_reg_1035_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1643
         assign bnn_RightShift_64Sx8S_1S_1_1643_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1643_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1644_in1 = {s_reg_1035_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1644
         assign bnn_RightShift_64Sx8S_1S_1_1644_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1644_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1645_in1 = {s_reg_1035_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1645
         assign bnn_RightShift_64Sx8S_1S_1_1645_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1645_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1646_in1 = {s_reg_1035_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1646
         assign bnn_RightShift_64Sx8S_1S_1_1646_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1646_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1647_in1 = {s_reg_1035_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1647
         assign bnn_RightShift_64Sx8S_1S_1_1647_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1647_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1648_in1 = {s_reg_1035_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1648
         assign bnn_RightShift_64Sx8S_1S_1_1648_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1648_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1649_in1 = {s_reg_1035_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1649
         assign bnn_RightShift_64Sx8S_1S_1_1649_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1649_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_4_1650_in1 = {s_reg_1035_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_1650
         assign bnn_RightShift_64Sx8S_1S_4_1650_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_1650_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1651_in1 = {s_reg_1039_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1651
         assign bnn_RightShift_64Sx8S_1S_1_1651_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1651_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1652_in1 = {s_reg_1039_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1652
         assign bnn_RightShift_64Sx8S_1S_1_1652_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1652_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1653_in1 = {s_reg_1039_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1653
         assign bnn_RightShift_64Sx8S_1S_1_1653_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1653_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1654_in1 = {s_reg_1039_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1654
         assign bnn_RightShift_64Sx8S_1S_1_1654_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1654_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1655_in1 = {s_reg_1039_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1655
         assign bnn_RightShift_64Sx8S_1S_1_1655_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1655_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1656_in1 = {s_reg_1039_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1656
         assign bnn_RightShift_64Sx8S_1S_1_1656_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1656_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1657_in1 = {s_reg_1039_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1657
         assign bnn_RightShift_64Sx8S_1S_1_1657_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1657_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1658_in1 = {s_reg_1039_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1658
         assign bnn_RightShift_64Sx8S_1S_1_1658_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1658_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1659_in1 = {s_reg_1027_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1659
         assign bnn_RightShift_64Sx8S_1S_1_1659_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1659_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1660_in1 = {s_reg_1027_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1660
         assign bnn_RightShift_64Sx8S_1S_1_1660_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1660_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1661_in1 = {s_reg_1027_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1661
         assign bnn_RightShift_64Sx8S_1S_1_1661_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1661_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1662_in1 = {s_reg_1027_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1662
         assign bnn_RightShift_64Sx8S_1S_1_1662_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1662_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1663_in1 = {s_reg_1027_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1663
         assign bnn_RightShift_64Sx8S_1S_1_1663_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1663_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1664_in1 = {s_reg_1027_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1664
         assign bnn_RightShift_64Sx8S_1S_1_1664_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1664_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1665_in1 = {s_reg_1027_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1665
         assign bnn_RightShift_64Sx8S_1S_1_1665_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1665_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1666_in1 = {s_reg_1027_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1666
         assign bnn_RightShift_64Sx8S_1S_1_1666_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1666_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1667_in1 = {s_reg_1047_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1667
         assign bnn_RightShift_64Sx8S_1S_1_1667_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1667_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1668_in1 = {s_reg_1047_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1668
         assign bnn_RightShift_64Sx8S_1S_1_1668_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1668_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1669_in1 = {s_reg_1047_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1669
         assign bnn_RightShift_64Sx8S_1S_1_1669_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1669_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1670_in1 = {s_reg_1047_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1670
         assign bnn_RightShift_64Sx8S_1S_1_1670_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1670_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1671_in1 = {s_reg_1047_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1671
         assign bnn_RightShift_64Sx8S_1S_1_1671_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1671_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1672_in1 = {s_reg_1047_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1672
         assign bnn_RightShift_64Sx8S_1S_1_1672_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1672_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1673_in1 = {s_reg_1047_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1673
         assign bnn_RightShift_64Sx8S_1S_1_1673_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1673_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_4_1674_in1 = {s_reg_1047_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_1674
         assign bnn_RightShift_64Sx8S_1S_4_1674_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_1674_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1675_in1 = {s_reg_1104[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1675
         assign bnn_RightShift_64Sx8S_1S_1_1675_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1675_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1676_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1675_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1676_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1676
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1676_out1_slice = bnn_N_Mux_3_2_6_1_1676_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1676_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1677
         assign bnn_RightShift_64Sx8S_1S_1_1677_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1103[5:0];

         assign bnn_N_Mux_3_2_6_1_1678_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1677_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1678_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1678
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1678_out1_slice = bnn_N_Mux_3_2_6_1_1678_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1678_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1679_in1 = {s_reg_1106[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1679
         assign bnn_RightShift_64Sx8S_1S_1_1679_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1679_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1680_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1679_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1680_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1680
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1680_out1_slice = bnn_N_Mux_3_2_6_1_1680_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1680_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1681
         assign bnn_RightShift_64Sx8S_1S_1_1681_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1105[5:0];

         assign bnn_N_Mux_3_2_6_1_1682_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1681_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1682_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1682
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1682_out1_slice = bnn_N_Mux_3_2_6_1_1682_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1682_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1683_in1 = {s_reg_1108, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1683
         assign bnn_RightShift_64Sx8S_1S_1_1683_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1683_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1684_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1683_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1684_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1684
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1684_out1_slice = bnn_N_Mux_3_2_6_1_1684_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1684_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1685
         assign bnn_RightShift_64Sx8S_1S_1_1685_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_Sub_8Sx2S_8S_4_1606_out1[5:0];

         assign bnn_N_Mux_3_2_6_1_1686_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1685_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1686_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1686
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1686_out1_slice = bnn_N_Mux_3_2_6_1_1686_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1686_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_1_1687_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[16], bnn_N_Mux_64_2_2_1_1636_out1[16]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1687_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1687
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1687_out1_slice = bnn_N_Mux_3_2_6_1_1687_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1687_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_3_2_6_1_1688_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[15], bnn_N_Mux_64_2_2_1_1636_out1[15]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1688_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1688
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1688_out1_slice = bnn_N_Mux_3_2_6_1_1688_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1688_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx7S_1S_1_1689_in1 = {s_reg_1070[3:0], 3'd0};

         // resource: bnn_RightShift_64Sx7S_1S_1  instance: bnn_RightShift_64Sx7S_1S_1_1689
         assign bnn_RightShift_64Sx7S_1S_1_1689_out1 = bnn_N_Mux_64_2_2_1_1636_out1 >> bnn_RightShift_64Sx7S_1S_1_1689_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1690_in1 = {s_reg_1070[4:0], 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1690
         assign bnn_RightShift_64Sx8S_1S_1_1690_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1690_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1691_in1 = {s_reg_1070[4:0], 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1691
         assign bnn_RightShift_64Sx8S_1S_1_1691_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1691_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1692_in1 = {s_reg_1070[4:0], 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1692
         assign bnn_RightShift_64Sx8S_1S_1_1692_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1692_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1693_in1 = {s_reg_1070[4:0], 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1693
         assign bnn_RightShift_64Sx8S_1S_1_1693_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1693_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1694_in1 = {s_reg_1070[4:0], 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1694
         assign bnn_RightShift_64Sx8S_1S_1_1694_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1694_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1695_in1 = {s_reg_1070[4:0], 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1695
         assign bnn_RightShift_64Sx8S_1S_1_1695_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1695_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1696_in1 = {s_reg_1070[4:0], 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1696
         assign bnn_RightShift_64Sx8S_1S_1_1696_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1696_in1[5:0];

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1697
         assign bnn_RightShift_64Sx8S_1S_1_1697_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1086[5:0];

         assign bnn_N_Mux_3_2_6_1_1698_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1697_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1698_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1698
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1698_out1_slice = bnn_N_Mux_3_2_6_1_1698_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1698_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1699_in1 = {s_reg_1036_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1699
         assign bnn_RightShift_64Sx8S_1S_1_1699_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1699_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1700_in1 = {s_reg_1036_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1700
         assign bnn_RightShift_64Sx8S_1S_1_1700_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1700_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1701_in1 = {s_reg_1036_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1701
         assign bnn_RightShift_64Sx8S_1S_1_1701_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1701_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1702_in1 = {s_reg_1036_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1702
         assign bnn_RightShift_64Sx8S_1S_1_1702_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1702_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1703_in1 = {s_reg_1036_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1703
         assign bnn_RightShift_64Sx8S_1S_1_1703_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1703_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1704_in1 = {s_reg_1036_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1704
         assign bnn_RightShift_64Sx8S_1S_1_1704_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1704_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1705_in1 = {s_reg_1036_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1705
         assign bnn_RightShift_64Sx8S_1S_1_1705_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1705_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1706_in1 = {s_reg_1036_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1706
         assign bnn_RightShift_64Sx8S_1S_1_1706_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1706_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1707_in1 = {s_reg_1030_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1707
         assign bnn_RightShift_64Sx8S_1S_1_1707_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1707_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1708_in1 = {s_reg_1030_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1708
         assign bnn_RightShift_64Sx8S_1S_1_1708_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1708_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1709_in1 = {s_reg_1030_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1709
         assign bnn_RightShift_64Sx8S_1S_1_1709_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1709_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1710_in1 = {s_reg_1030_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1710
         assign bnn_RightShift_64Sx8S_1S_1_1710_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1710_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1711_in1 = {s_reg_1030_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1711
         assign bnn_RightShift_64Sx8S_1S_1_1711_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1711_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1712_in1 = {s_reg_1030_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1712
         assign bnn_RightShift_64Sx8S_1S_1_1712_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1712_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1713_in1 = {s_reg_1030_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1713
         assign bnn_RightShift_64Sx8S_1S_1_1713_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1713_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1714_in1 = {s_reg_1030_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1714
         assign bnn_RightShift_64Sx8S_1S_1_1714_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1714_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1715_in1 = {s_reg_1043_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1715
         assign bnn_RightShift_64Sx8S_1S_1_1715_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1715_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1716_in1 = {s_reg_1043_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1716
         assign bnn_RightShift_64Sx8S_1S_1_1716_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1716_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1717_in1 = {s_reg_1043_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1717
         assign bnn_RightShift_64Sx8S_1S_1_1717_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1717_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1718_in1 = {s_reg_1043_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1718
         assign bnn_RightShift_64Sx8S_1S_1_1718_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1718_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1719_in1 = {s_reg_1043_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1719
         assign bnn_RightShift_64Sx8S_1S_1_1719_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1719_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1720_in1 = {s_reg_1043_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1720
         assign bnn_RightShift_64Sx8S_1S_1_1720_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1720_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1721_in1 = {s_reg_1043_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1721
         assign bnn_RightShift_64Sx8S_1S_1_1721_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1721_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1722_in1 = {s_reg_1043_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1722
         assign bnn_RightShift_64Sx8S_1S_1_1722_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1722_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1723_in1 = {s_reg_871_stage1, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1723
         assign bnn_RightShift_64Sx8S_1S_1_1723_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1723_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1724_in1 = {s_reg_871_stage1, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1724
         assign bnn_RightShift_64Sx8S_1S_1_1724_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1724_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1725_in1 = {s_reg_871_stage1, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1725
         assign bnn_RightShift_64Sx8S_1S_1_1725_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1725_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1726_in1 = {s_reg_871_stage1, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1726
         assign bnn_RightShift_64Sx8S_1S_1_1726_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1726_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1727_in1 = {s_reg_871_stage1, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1727
         assign bnn_RightShift_64Sx8S_1S_1_1727_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1727_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1728_in1 = {s_reg_871_stage1, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1728
         assign bnn_RightShift_64Sx8S_1S_1_1728_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1728_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1729_in1 = {s_reg_871_stage1, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1729
         assign bnn_RightShift_64Sx8S_1S_1_1729_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1729_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_4_1730_in1 = {s_reg_871_stage1, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_1730
         assign bnn_RightShift_64Sx8S_1S_4_1730_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_1730_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1731_in1 = {s_reg_1021_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1731
         assign bnn_RightShift_64Sx8S_1S_1_1731_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1731_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1732_in1 = {s_reg_1021_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1732
         assign bnn_RightShift_64Sx8S_1S_1_1732_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1732_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1733_in1 = {s_reg_1021_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1733
         assign bnn_RightShift_64Sx8S_1S_1_1733_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1733_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1734_in1 = {s_reg_1021_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1734
         assign bnn_RightShift_64Sx8S_1S_1_1734_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1734_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1735_in1 = {s_reg_1021_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1735
         assign bnn_RightShift_64Sx8S_1S_1_1735_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1735_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1736_in1 = {s_reg_1021_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1736
         assign bnn_RightShift_64Sx8S_1S_1_1736_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1736_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1737_in1 = {s_reg_1021_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1737
         assign bnn_RightShift_64Sx8S_1S_1_1737_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1737_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1738_in1 = {s_reg_1021_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1738
         assign bnn_RightShift_64Sx8S_1S_1_1738_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1738_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1739_in1 = {s_reg_1031_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1739
         assign bnn_RightShift_64Sx8S_1S_1_1739_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1739_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1740_in1 = {s_reg_1031_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1740
         assign bnn_RightShift_64Sx8S_1S_1_1740_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1740_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1741_in1 = {s_reg_1031_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1741
         assign bnn_RightShift_64Sx8S_1S_1_1741_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1741_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1742_in1 = {s_reg_1031_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1742
         assign bnn_RightShift_64Sx8S_1S_1_1742_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1742_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1743_in1 = {s_reg_1031_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1743
         assign bnn_RightShift_64Sx8S_1S_1_1743_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1743_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1744_in1 = {s_reg_1031_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1744
         assign bnn_RightShift_64Sx8S_1S_1_1744_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1744_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1745_in1 = {s_reg_1031_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1745
         assign bnn_RightShift_64Sx8S_1S_1_1745_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1745_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1746_in1 = {s_reg_1031_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1746
         assign bnn_RightShift_64Sx8S_1S_1_1746_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1746_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1747_in1 = {s_reg_1046_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1747
         assign bnn_RightShift_64Sx8S_1S_1_1747_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1747_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1748_in1 = {s_reg_1046_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1748
         assign bnn_RightShift_64Sx8S_1S_1_1748_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1748_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1749_in1 = {s_reg_1046_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1749
         assign bnn_RightShift_64Sx8S_1S_1_1749_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1749_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1750_in1 = {s_reg_1046_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1750
         assign bnn_RightShift_64Sx8S_1S_1_1750_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1750_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1751_in1 = {s_reg_1046_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1751
         assign bnn_RightShift_64Sx8S_1S_1_1751_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1751_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1752_in1 = {s_reg_1046_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1752
         assign bnn_RightShift_64Sx8S_1S_1_1752_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1752_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1753_in1 = {s_reg_1046_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1753
         assign bnn_RightShift_64Sx8S_1S_1_1753_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1753_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_4_1754_in1 = {s_reg_1046_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_1754
         assign bnn_RightShift_64Sx8S_1S_4_1754_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_1754_in1[5:0];

         assign bnn_RightShift_64Sx8S_1S_1_1755_in1 = {s_reg_874[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1755
         assign bnn_RightShift_64Sx8S_1S_1_1755_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1755_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1756_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1755_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1756_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1756
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1756_out1_slice = bnn_N_Mux_3_2_6_1_1756_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1756_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1757_in1 = {s_reg_1091[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1757
         assign bnn_RightShift_64Sx8S_1S_1_1757_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1757_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1758_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1757_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1758_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1758
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1758_out1_slice = bnn_N_Mux_3_2_6_1_1758_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1758_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1759
         assign bnn_RightShift_64Sx8S_1S_1_1759_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1090[5:0];

         assign bnn_N_Mux_3_2_6_1_1760_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1759_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1760_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1760
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1760_out1_slice = bnn_N_Mux_3_2_6_1_1760_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1760_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1761_in1 = {s_reg_1099, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1761
         assign bnn_RightShift_64Sx8S_1S_1_1761_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1761_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1762_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1761_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1762_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1762
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1762_out1_slice = bnn_N_Mux_3_2_6_1_1762_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1762_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1763
         assign bnn_RightShift_64Sx8S_1S_1_1763_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1098[5:0];

         assign bnn_N_Mux_3_2_6_1_1764_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1763_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1764_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1764
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1764_out1_slice = bnn_N_Mux_3_2_6_1_1764_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1764_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1765_in1 = {s_reg_1095[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1765
         assign bnn_RightShift_64Sx8S_1S_1_1765_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1765_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1766_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1765_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1766_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1766
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1766_out1_slice = bnn_N_Mux_3_2_6_1_1766_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1766_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1767
         assign bnn_RightShift_64Sx8S_1S_1_1767_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1092[5:0];

         assign bnn_N_Mux_3_2_6_1_1768_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1767_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1768_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1768
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1768_out1_slice = bnn_N_Mux_3_2_6_1_1768_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1768_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1769_in1 = {s_reg_1101[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1769
         assign bnn_RightShift_64Sx8S_1S_1_1769_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1769_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1770_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1769_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1770_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1770
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1770_out1_slice = bnn_N_Mux_3_2_6_1_1770_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1770_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1771
         assign bnn_RightShift_64Sx8S_1S_1_1771_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1100[5:0];

         assign bnn_N_Mux_3_2_6_1_1772_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1771_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_1772_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_1772
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_1772_out1_slice = bnn_N_Mux_3_2_6_1_1772_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1772_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1773_in1 = {s_reg_1102[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1773
         assign bnn_RightShift_64Sx8S_1S_1_1773_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1773_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_1774_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1773_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1774_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1774
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1774_out1_slice = bnn_N_Mux_3_2_6_1_1774_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1774_out1_slice = 2'd0;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1775
         assign bnn_RightShift_64Sx8S_1S_1_1775_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_Sub_8Sx2S_8S_4_1596_out1[5:0];

         assign bnn_N_Mux_3_2_6_1_1776_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1775_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1776_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1776
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1776_out1_slice = bnn_N_Mux_3_2_6_1_1776_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1776_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1777_in1 = {s_reg_1068_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1777
         assign bnn_RightShift_64Sx8S_1S_1_1777_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1777_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1778_in3 = {bnn_RightShift_64Sx8S_1S_1_1777_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_872 or bnn_N_Mux_2_2_3_1_1778_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1778
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1778_out1 = s_reg_872;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1778_out1 = bnn_N_Mux_2_2_3_1_1778_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_874[1:0] or s_reg_876 or s_reg_879 or bnn_N_Mux_2_2_3_1_1778_out1)
          begin :bnn_N_Mux_2_4_8_1_1779
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1779_out1 = bnn_N_Mux_2_2_3_1_1778_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1779_out1 = s_reg_876;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1779_out1 = s_reg_874[1:0];
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1779_out1 = s_reg_879;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1779_out1)
          begin :bnn_N_Mux_3_2_6_1_1780
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1780_out1_slice = bnn_N_Mux_2_4_8_1_1779_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1780_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1781_in3 = {bnn_RightShift_64Sx7S_1S_1_1689_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1781_in3 or bnn_N_Mux_3_2_6_1_1780_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1781
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1781_out1 = bnn_N_Mux_3_2_6_1_1780_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1781_out1 = bnn_N_Mux_2_2_3_1_1781_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_9_4
         always @(s_reg_1004 or s_reg_977 or s_reg_984 or bnn_N_Mux_2_2_3_1_1781_out1)
          begin :bnn_N_Mux_2_4_9_4_1782
            case (s_reg_1004) 

               2'd0: begin
                  bnn_N_Mux_2_4_9_4_1782_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_9_4_1782_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_9_4_1782_out1 = s_reg_984;
               end
               
               default: begin
                  bnn_N_Mux_2_4_9_4_1782_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_And_1Sx1U_1U_4_1584_out1 or bnn_N_Mux_2_4_9_4_1782_out1)
          begin :bnn_N_Mux_3_2_6_1_1783
            if (bnn_And_1Sx1U_1U_4_1584_out1) begin
               bnn_N_Mux_3_2_6_1_1783_out1_slice = bnn_N_Mux_2_4_9_4_1782_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1783_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_9_4
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_1781_out1 or bnn_N_Mux_3_2_6_1_1783_out1_slice)
          begin :bnn_N_Mux_2_4_9_4_1784
            case (s_reg_1004) 

               2'd0: begin
                  bnn_N_Mux_2_4_9_4_1784_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_9_4_1784_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_9_4_1784_out1 = bnn_N_Mux_3_2_6_1_1783_out1_slice;
               end
               
               default: begin
                  bnn_N_Mux_2_4_9_4_1784_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_And_1Sx1U_1U_4_1585_out1 or bnn_N_Mux_2_4_9_4_1784_out1)
          begin :bnn_N_Mux_3_2_6_1_1785
            if (bnn_And_1Sx1U_1U_4_1585_out1) begin
               bnn_N_Mux_3_2_6_1_1785_out1_slice = bnn_N_Mux_2_4_9_4_1784_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1785_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1786_in1 = {s_reg_1068_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1786
         assign bnn_RightShift_64Sx8S_1S_1_1786_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1786_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1787_in3 = {bnn_RightShift_64Sx8S_1S_1_1786_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_873 or bnn_N_Mux_2_2_3_1_1787_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1787
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1787_out1 = s_reg_873;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1787_out1 = bnn_N_Mux_2_2_3_1_1787_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_875 or s_reg_877 or s_reg_880 or bnn_N_Mux_2_2_3_1_1787_out1)
          begin :bnn_N_Mux_2_4_8_1_1788
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1788_out1 = bnn_N_Mux_2_2_3_1_1787_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1788_out1 = s_reg_877;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1788_out1 = s_reg_875;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1788_out1 = s_reg_880;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1788_out1)
          begin :bnn_N_Mux_3_2_6_1_1789
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1789_out1_slice = bnn_N_Mux_2_4_8_1_1788_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1789_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1790_in3 = {bnn_RightShift_64Sx8S_1S_1_1690_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1790_in3 or bnn_N_Mux_3_2_6_1_1789_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1790
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1790_out1 = bnn_N_Mux_3_2_6_1_1789_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1790_out1 = bnn_N_Mux_2_2_3_1_1790_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1791_in1 = {s_reg_1068_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1791
         assign bnn_RightShift_64Sx8S_1S_1_1791_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1791_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1792_in3 = {bnn_RightShift_64Sx8S_1S_1_1791_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_878 or bnn_N_Mux_2_2_3_1_1792_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1792
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1792_out1 = s_reg_878;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1792_out1 = bnn_N_Mux_2_2_3_1_1792_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_881 or s_reg_882 or s_reg_885 or bnn_N_Mux_2_2_3_1_1792_out1)
          begin :bnn_N_Mux_2_4_8_1_1793
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1793_out1 = bnn_N_Mux_2_2_3_1_1792_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1793_out1 = s_reg_882;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1793_out1 = s_reg_881;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1793_out1 = s_reg_885;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1793_out1)
          begin :bnn_N_Mux_3_2_6_1_1794
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1794_out1_slice = bnn_N_Mux_2_4_8_1_1793_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1794_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1795_in3 = {bnn_RightShift_64Sx8S_1S_1_1691_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1795_in3 or bnn_N_Mux_3_2_6_1_1794_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1795
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1795_out1 = bnn_N_Mux_3_2_6_1_1794_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1795_out1 = bnn_N_Mux_2_2_3_1_1795_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1796_in1 = {s_reg_1068_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1796
         assign bnn_RightShift_64Sx8S_1S_1_1796_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1796_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1797_in3 = {bnn_RightShift_64Sx8S_1S_1_1796_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_884 or bnn_N_Mux_2_2_3_1_1797_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1797
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1797_out1 = s_reg_884;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1797_out1 = bnn_N_Mux_2_2_3_1_1797_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_888 or s_reg_889 or s_reg_892 or bnn_N_Mux_2_2_3_1_1797_out1)
          begin :bnn_N_Mux_2_4_8_1_1798
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1798_out1 = bnn_N_Mux_2_2_3_1_1797_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1798_out1 = s_reg_889;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1798_out1 = s_reg_888;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1798_out1 = s_reg_892;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1798_out1)
          begin :bnn_N_Mux_3_2_6_1_1799
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1799_out1_slice = bnn_N_Mux_2_4_8_1_1798_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1799_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1800_in3 = {bnn_RightShift_64Sx8S_1S_1_1692_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1800_in3 or bnn_N_Mux_3_2_6_1_1799_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1800
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1800_out1 = bnn_N_Mux_3_2_6_1_1799_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1800_out1 = bnn_N_Mux_2_2_3_1_1800_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1801_in1 = {s_reg_1068_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1801
         assign bnn_RightShift_64Sx8S_1S_1_1801_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1801_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1802_in3 = {bnn_RightShift_64Sx8S_1S_1_1801_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_890 or bnn_N_Mux_2_2_3_1_1802_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1802
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1802_out1 = s_reg_890;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1802_out1 = bnn_N_Mux_2_2_3_1_1802_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_898 or s_reg_899 or s_reg_901 or bnn_N_Mux_2_2_3_1_1802_out1)
          begin :bnn_N_Mux_2_4_8_1_1803
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1803_out1 = bnn_N_Mux_2_2_3_1_1802_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1803_out1 = s_reg_899;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1803_out1 = s_reg_898;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1803_out1 = s_reg_901;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1803_out1)
          begin :bnn_N_Mux_3_2_6_1_1804
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1804_out1_slice = bnn_N_Mux_2_4_8_1_1803_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1804_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1805_in3 = {bnn_RightShift_64Sx8S_1S_1_1693_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1805_in3 or bnn_N_Mux_3_2_6_1_1804_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1805
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1805_out1 = bnn_N_Mux_3_2_6_1_1804_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1805_out1 = bnn_N_Mux_2_2_3_1_1805_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1806_in1 = {s_reg_1068_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1806
         assign bnn_RightShift_64Sx8S_1S_1_1806_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1806_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1807_in3 = {bnn_RightShift_64Sx8S_1S_1_1806_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_900 or bnn_N_Mux_2_2_3_1_1807_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1807
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1807_out1 = s_reg_900;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1807_out1 = bnn_N_Mux_2_2_3_1_1807_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_909 or s_reg_910 or s_reg_912 or bnn_N_Mux_2_2_3_1_1807_out1)
          begin :bnn_N_Mux_2_4_8_1_1808
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1808_out1 = bnn_N_Mux_2_2_3_1_1807_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1808_out1 = s_reg_910;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1808_out1 = s_reg_909;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1808_out1 = s_reg_912;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1808_out1)
          begin :bnn_N_Mux_3_2_6_1_1809
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1809_out1_slice = bnn_N_Mux_2_4_8_1_1808_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1809_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1810_in3 = {bnn_RightShift_64Sx8S_1S_1_1694_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1810_in3 or bnn_N_Mux_3_2_6_1_1809_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1810
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1810_out1 = bnn_N_Mux_3_2_6_1_1809_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1810_out1 = bnn_N_Mux_2_2_3_1_1810_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1811_in1 = {s_reg_1068_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1811
         assign bnn_RightShift_64Sx8S_1S_1_1811_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1811_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1812_in3 = {bnn_RightShift_64Sx8S_1S_1_1811_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_911 or bnn_N_Mux_2_2_3_1_1812_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1812
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1812_out1 = s_reg_911;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1812_out1 = bnn_N_Mux_2_2_3_1_1812_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_917 or s_reg_918 or s_reg_920 or bnn_N_Mux_2_2_3_1_1812_out1)
          begin :bnn_N_Mux_2_4_8_1_1813
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1813_out1 = bnn_N_Mux_2_2_3_1_1812_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1813_out1 = s_reg_918;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1813_out1 = s_reg_917;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1813_out1 = s_reg_920;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1813_out1)
          begin :bnn_N_Mux_3_2_6_1_1814
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1814_out1_slice = bnn_N_Mux_2_4_8_1_1813_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1814_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1815_in3 = {bnn_RightShift_64Sx8S_1S_1_1695_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1815_in3 or bnn_N_Mux_3_2_6_1_1814_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1815
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1815_out1 = bnn_N_Mux_3_2_6_1_1814_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1815_out1 = bnn_N_Mux_2_2_3_1_1815_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1816_in1 = {s_reg_1068_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1816
         assign bnn_RightShift_64Sx8S_1S_1_1816_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1816_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1817_in3 = {bnn_RightShift_64Sx8S_1S_1_1816_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_919 or bnn_N_Mux_2_2_3_1_1817_in3 or s_reg_1069_stage1)
          begin :bnn_N_Mux_2_2_3_1_1817
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_1817_out1 = s_reg_919;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1817_out1 = bnn_N_Mux_2_2_3_1_1817_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_925 or s_reg_926 or s_reg_928 or bnn_N_Mux_2_2_3_1_1817_out1)
          begin :bnn_N_Mux_2_4_8_1_1818
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1818_out1 = bnn_N_Mux_2_2_3_1_1817_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1818_out1 = s_reg_926;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1818_out1 = s_reg_925;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1818_out1 = s_reg_928;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_1818_out1)
          begin :bnn_N_Mux_3_2_6_1_1819
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_1819_out1_slice = bnn_N_Mux_2_4_8_1_1818_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_1819_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1820_in3 = {bnn_RightShift_64Sx8S_1S_1_1696_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_2_2_3_1_1820_in3 or bnn_N_Mux_3_2_6_1_1819_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1820
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_1820_out1 = bnn_N_Mux_3_2_6_1_1819_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1820_out1 = bnn_N_Mux_2_2_3_1_1820_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1821_in1 = {s_reg_1076_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1821
         assign bnn_RightShift_64Sx8S_1S_1_1821_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1821_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1822_in3 = {bnn_RightShift_64Sx8S_1S_1_1821_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_886[1:0] or bnn_N_Mux_2_2_3_1_1822_in3)
          begin :bnn_N_Mux_2_2_3_1_1822
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1822_out1 = s_reg_886[1:0];
            end
            else begin
               bnn_N_Mux_2_2_3_1_1822_out1 = bnn_N_Mux_2_2_3_1_1822_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_879 or s_reg_893 or s_reg_896 or bnn_N_Mux_2_2_3_1_1822_out1)
          begin :bnn_N_Mux_2_4_8_1_1823
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1823_out1 = bnn_N_Mux_2_2_3_1_1822_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1823_out1 = s_reg_893;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1823_out1 = s_reg_879;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1823_out1 = s_reg_896;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1823_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1824
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1824_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1824_out1 = bnn_N_Mux_2_4_8_1_1823_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1825_in3 = {bnn_RightShift_64Sx8S_1S_1_1699_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1824_out1 or bnn_N_Mux_2_2_3_1_1825_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1825
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1825_out1 = bnn_N_Mux_2_2_3_1_1824_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1825_out1 = bnn_N_Mux_2_2_3_1_1825_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1826_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[0], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1778_out1 or bnn_N_Mux_2_2_3_1_1781_out1 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_N_Mux_2_4_8_1_1826_in3)
          begin :bnn_N_Mux_2_4_8_1_1826
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1826_out1 = bnn_N_Mux_2_2_3_1_1778_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1826_out1 = bnn_N_Mux_2_4_8_1_1826_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1826_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1826_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1826_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1827
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1827_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1827_out1 = bnn_N_Mux_2_4_8_1_1826_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1828_in3 = {bnn_RightShift_64Sx8S_1S_1_1723_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1827_out1 or bnn_N_Mux_2_2_3_1_1828_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1828
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1828_out1 = bnn_N_Mux_2_2_3_1_1827_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1828_out1 = bnn_N_Mux_2_2_3_1_1828_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1781_out1 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_N_Mux_2_4_8_1_1826_in3 or bnn_N_Mux_2_2_3_1_1828_out1)
          begin :bnn_N_Mux_2_4_8_1_1829
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1829_out1 = bnn_N_Mux_2_2_3_1_1828_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1829_out1 = bnn_N_Mux_2_4_8_1_1826_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1829_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1829_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1829_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1830
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1830_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1830_out1 = bnn_N_Mux_2_4_8_1_1829_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1831_in3 = {bnn_RightShift_64Sx8S_1S_1_1643_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1830_out1 or bnn_N_Mux_2_2_3_1_1831_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1831
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1831_out1 = bnn_N_Mux_2_2_3_1_1830_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1831_out1 = bnn_N_Mux_2_2_3_1_1831_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_9_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1831_out1 or bnn_N_Mux_3_2_6_1_1783_out1_slice or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_9_4_1832
            case (s_reg_1004) 

               2'd0: begin
                  bnn_N_Mux_2_4_9_4_1832_out1 = bnn_N_Mux_2_2_3_1_1831_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_9_4_1832_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_9_4_1832_out1 = bnn_N_Mux_3_2_6_1_1783_out1_slice;
               end
               
               default: begin
                  bnn_N_Mux_2_4_9_4_1832_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_1587_out1 or bnn_N_Mux_2_4_9_4_1832_out1)
          begin :bnn_N_Mux_3_2_6_4_1833
            if (bnn_And_1Sx1U_1U_4_1587_out1) begin
               bnn_N_Mux_3_2_6_4_1833_out1_slice = bnn_N_Mux_2_4_9_4_1832_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_1833_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_9_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1831_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice or bnn_N_Mux_3_2_6_4_1833_out1_slice)
          begin :bnn_N_Mux_2_4_9_4_1834
            case (s_reg_1004) 

               2'd0: begin
                  bnn_N_Mux_2_4_9_4_1834_out1 = bnn_N_Mux_2_2_3_1_1831_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_9_4_1834_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_9_4_1834_out1 = bnn_N_Mux_3_2_6_4_1833_out1_slice;
               end
               
               default: begin
                  bnn_N_Mux_2_4_9_4_1834_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_1630_out1 or bnn_N_Mux_2_4_9_4_1834_out1)
          begin :bnn_N_Mux_3_2_6_4_1835
            if (bnn_And_1Sx1U_1U_4_1630_out1) begin
               bnn_N_Mux_3_2_6_4_1835_out1_slice = bnn_N_Mux_2_4_9_4_1834_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_1835_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1836_in1 = {s_reg_1076_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1836
         assign bnn_RightShift_64Sx8S_1S_1_1836_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1836_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1837_in3 = {bnn_RightShift_64Sx8S_1S_1_1836_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_895 or bnn_N_Mux_2_2_3_1_1837_in3)
          begin :bnn_N_Mux_2_2_3_1_1837
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1837_out1 = s_reg_895;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1837_out1 = bnn_N_Mux_2_2_3_1_1837_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_880 or s_reg_903 or s_reg_906 or bnn_N_Mux_2_2_3_1_1837_out1)
          begin :bnn_N_Mux_2_4_8_1_1838
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1838_out1 = bnn_N_Mux_2_2_3_1_1837_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1838_out1 = s_reg_903;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1838_out1 = s_reg_880;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1838_out1 = s_reg_906;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1838_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1839
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1839_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1839_out1 = bnn_N_Mux_2_4_8_1_1838_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1840_in3 = {bnn_RightShift_64Sx8S_1S_1_1700_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1839_out1 or bnn_N_Mux_2_2_3_1_1840_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1840
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1840_out1 = bnn_N_Mux_2_2_3_1_1839_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1840_out1 = bnn_N_Mux_2_2_3_1_1840_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1841_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[1], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1787_out1 or bnn_N_Mux_2_2_3_1_1790_out1 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_N_Mux_2_4_8_1_1841_in3)
          begin :bnn_N_Mux_2_4_8_1_1841
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1841_out1 = bnn_N_Mux_2_2_3_1_1787_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1841_out1 = bnn_N_Mux_2_4_8_1_1841_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1841_out1 = bnn_N_Mux_2_2_3_1_1790_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1841_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1841_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1842
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1842_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1842_out1 = bnn_N_Mux_2_4_8_1_1841_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1843_in3 = {bnn_RightShift_64Sx8S_1S_1_1724_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1842_out1 or bnn_N_Mux_2_2_3_1_1843_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1843
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1843_out1 = bnn_N_Mux_2_2_3_1_1842_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1843_out1 = bnn_N_Mux_2_2_3_1_1843_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1790_out1 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_N_Mux_2_4_8_1_1841_in3 or bnn_N_Mux_2_2_3_1_1843_out1)
          begin :bnn_N_Mux_2_4_8_1_1844
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1844_out1 = bnn_N_Mux_2_2_3_1_1843_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1844_out1 = bnn_N_Mux_2_4_8_1_1841_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1844_out1 = bnn_N_Mux_2_2_3_1_1790_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1844_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1844_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1845
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1845_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1845_out1 = bnn_N_Mux_2_4_8_1_1844_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1846_in3 = {bnn_RightShift_64Sx8S_1S_1_1644_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1845_out1 or bnn_N_Mux_2_2_3_1_1846_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1846
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1846_out1 = bnn_N_Mux_2_2_3_1_1845_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1846_out1 = bnn_N_Mux_2_2_3_1_1846_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1847_in1 = {s_reg_1076_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1847
         assign bnn_RightShift_64Sx8S_1S_1_1847_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1847_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1848_in3 = {bnn_RightShift_64Sx8S_1S_1_1847_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_904 or bnn_N_Mux_2_2_3_1_1848_in3)
          begin :bnn_N_Mux_2_2_3_1_1848
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1848_out1 = s_reg_904;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1848_out1 = bnn_N_Mux_2_2_3_1_1848_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_885 or s_reg_913 or s_reg_915 or bnn_N_Mux_2_2_3_1_1848_out1)
          begin :bnn_N_Mux_2_4_8_1_1849
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1849_out1 = bnn_N_Mux_2_2_3_1_1848_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1849_out1 = s_reg_913;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1849_out1 = s_reg_885;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1849_out1 = s_reg_915;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1849_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1850
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1850_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1850_out1 = bnn_N_Mux_2_4_8_1_1849_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1851_in3 = {bnn_RightShift_64Sx8S_1S_1_1701_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1850_out1 or bnn_N_Mux_2_2_3_1_1851_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1851
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1851_out1 = bnn_N_Mux_2_2_3_1_1850_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1851_out1 = bnn_N_Mux_2_2_3_1_1851_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1852_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[2], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1792_out1 or bnn_N_Mux_2_2_3_1_1795_out1 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_N_Mux_2_4_8_1_1852_in3)
          begin :bnn_N_Mux_2_4_8_1_1852
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1852_out1 = bnn_N_Mux_2_2_3_1_1792_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1852_out1 = bnn_N_Mux_2_4_8_1_1852_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1852_out1 = bnn_N_Mux_2_2_3_1_1795_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1852_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1852_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1853
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1853_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1853_out1 = bnn_N_Mux_2_4_8_1_1852_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1854_in3 = {bnn_RightShift_64Sx8S_1S_1_1725_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1853_out1 or bnn_N_Mux_2_2_3_1_1854_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1854
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1854_out1 = bnn_N_Mux_2_2_3_1_1853_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1854_out1 = bnn_N_Mux_2_2_3_1_1854_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1795_out1 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_N_Mux_2_4_8_1_1852_in3 or bnn_N_Mux_2_2_3_1_1854_out1)
          begin :bnn_N_Mux_2_4_8_1_1855
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1855_out1 = bnn_N_Mux_2_2_3_1_1854_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1855_out1 = bnn_N_Mux_2_4_8_1_1852_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1855_out1 = bnn_N_Mux_2_2_3_1_1795_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1855_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1855_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1856
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1856_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1856_out1 = bnn_N_Mux_2_4_8_1_1855_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1857_in3 = {bnn_RightShift_64Sx8S_1S_1_1645_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1856_out1 or bnn_N_Mux_2_2_3_1_1857_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1857
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1857_out1 = bnn_N_Mux_2_2_3_1_1856_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1857_out1 = bnn_N_Mux_2_2_3_1_1857_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1858_in1 = {s_reg_1076_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1858
         assign bnn_RightShift_64Sx8S_1S_1_1858_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1858_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1859_in3 = {bnn_RightShift_64Sx8S_1S_1_1858_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_914 or bnn_N_Mux_2_2_3_1_1859_in3)
          begin :bnn_N_Mux_2_2_3_1_1859
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1859_out1 = s_reg_914;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1859_out1 = bnn_N_Mux_2_2_3_1_1859_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_892 or s_reg_921 or s_reg_923 or bnn_N_Mux_2_2_3_1_1859_out1)
          begin :bnn_N_Mux_2_4_8_1_1860
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1860_out1 = bnn_N_Mux_2_2_3_1_1859_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1860_out1 = s_reg_921;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1860_out1 = s_reg_892;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1860_out1 = s_reg_923;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1860_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1861
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1861_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1861_out1 = bnn_N_Mux_2_4_8_1_1860_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1862_in3 = {bnn_RightShift_64Sx8S_1S_1_1702_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1861_out1 or bnn_N_Mux_2_2_3_1_1862_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1862
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1862_out1 = bnn_N_Mux_2_2_3_1_1861_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1862_out1 = bnn_N_Mux_2_2_3_1_1862_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1863_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[3], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1797_out1 or bnn_N_Mux_2_2_3_1_1800_out1 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_N_Mux_2_4_8_1_1863_in3)
          begin :bnn_N_Mux_2_4_8_1_1863
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1863_out1 = bnn_N_Mux_2_2_3_1_1797_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1863_out1 = bnn_N_Mux_2_4_8_1_1863_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1863_out1 = bnn_N_Mux_2_2_3_1_1800_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1863_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1863_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1864
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1864_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1864_out1 = bnn_N_Mux_2_4_8_1_1863_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1865_in3 = {bnn_RightShift_64Sx8S_1S_1_1726_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1864_out1 or bnn_N_Mux_2_2_3_1_1865_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1865
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1865_out1 = bnn_N_Mux_2_2_3_1_1864_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1865_out1 = bnn_N_Mux_2_2_3_1_1865_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1800_out1 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_N_Mux_2_4_8_1_1863_in3 or bnn_N_Mux_2_2_3_1_1865_out1)
          begin :bnn_N_Mux_2_4_8_1_1866
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1866_out1 = bnn_N_Mux_2_2_3_1_1865_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1866_out1 = bnn_N_Mux_2_4_8_1_1863_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1866_out1 = bnn_N_Mux_2_2_3_1_1800_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1866_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1866_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1867
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1867_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1867_out1 = bnn_N_Mux_2_4_8_1_1866_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1868_in3 = {bnn_RightShift_64Sx8S_1S_1_1646_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1867_out1 or bnn_N_Mux_2_2_3_1_1868_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1868
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1868_out1 = bnn_N_Mux_2_2_3_1_1867_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1868_out1 = bnn_N_Mux_2_2_3_1_1868_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1869_in1 = {s_reg_1076_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1869
         assign bnn_RightShift_64Sx8S_1S_1_1869_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1869_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1870_in3 = {bnn_RightShift_64Sx8S_1S_1_1869_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_922 or bnn_N_Mux_2_2_3_1_1870_in3)
          begin :bnn_N_Mux_2_2_3_1_1870
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1870_out1 = s_reg_922;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1870_out1 = bnn_N_Mux_2_2_3_1_1870_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_901 or s_reg_929 or s_reg_931 or bnn_N_Mux_2_2_3_1_1870_out1)
          begin :bnn_N_Mux_2_4_8_1_1871
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1871_out1 = bnn_N_Mux_2_2_3_1_1870_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1871_out1 = s_reg_929;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1871_out1 = s_reg_901;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1871_out1 = s_reg_931;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1871_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1872
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1872_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1872_out1 = bnn_N_Mux_2_4_8_1_1871_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1873_in3 = {bnn_RightShift_64Sx8S_1S_1_1703_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1872_out1 or bnn_N_Mux_2_2_3_1_1873_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1873
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1873_out1 = bnn_N_Mux_2_2_3_1_1872_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1873_out1 = bnn_N_Mux_2_2_3_1_1873_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1874_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[4], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1802_out1 or bnn_N_Mux_2_2_3_1_1805_out1 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_N_Mux_2_4_8_1_1874_in3)
          begin :bnn_N_Mux_2_4_8_1_1874
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1874_out1 = bnn_N_Mux_2_2_3_1_1802_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1874_out1 = bnn_N_Mux_2_4_8_1_1874_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1874_out1 = bnn_N_Mux_2_2_3_1_1805_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1874_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1874_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1875
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1875_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1875_out1 = bnn_N_Mux_2_4_8_1_1874_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1876_in3 = {bnn_RightShift_64Sx8S_1S_1_1727_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1875_out1 or bnn_N_Mux_2_2_3_1_1876_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1876
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1876_out1 = bnn_N_Mux_2_2_3_1_1875_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1876_out1 = bnn_N_Mux_2_2_3_1_1876_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1805_out1 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_N_Mux_2_4_8_1_1874_in3 or bnn_N_Mux_2_2_3_1_1876_out1)
          begin :bnn_N_Mux_2_4_8_1_1877
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1877_out1 = bnn_N_Mux_2_2_3_1_1876_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1877_out1 = bnn_N_Mux_2_4_8_1_1874_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1877_out1 = bnn_N_Mux_2_2_3_1_1805_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1877_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1877_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1878
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1878_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1878_out1 = bnn_N_Mux_2_4_8_1_1877_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1879_in3 = {bnn_RightShift_64Sx8S_1S_1_1647_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1878_out1 or bnn_N_Mux_2_2_3_1_1879_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1879
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1879_out1 = bnn_N_Mux_2_2_3_1_1878_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1879_out1 = bnn_N_Mux_2_2_3_1_1879_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1880_in1 = {s_reg_1076_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1880
         assign bnn_RightShift_64Sx8S_1S_1_1880_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1880_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1881_in3 = {bnn_RightShift_64Sx8S_1S_1_1880_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_930 or bnn_N_Mux_2_2_3_1_1881_in3)
          begin :bnn_N_Mux_2_2_3_1_1881
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1881_out1 = s_reg_930;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1881_out1 = bnn_N_Mux_2_2_3_1_1881_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_912 or s_reg_936 or s_reg_938 or bnn_N_Mux_2_2_3_1_1881_out1)
          begin :bnn_N_Mux_2_4_8_1_1882
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1882_out1 = bnn_N_Mux_2_2_3_1_1881_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1882_out1 = s_reg_936;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1882_out1 = s_reg_912;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1882_out1 = s_reg_938;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1882_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1883
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1883_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1883_out1 = bnn_N_Mux_2_4_8_1_1882_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1884_in3 = {bnn_RightShift_64Sx8S_1S_1_1704_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1883_out1 or bnn_N_Mux_2_2_3_1_1884_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1884
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1884_out1 = bnn_N_Mux_2_2_3_1_1883_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1884_out1 = bnn_N_Mux_2_2_3_1_1884_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1885_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[5], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1807_out1 or bnn_N_Mux_2_2_3_1_1810_out1 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_N_Mux_2_4_8_1_1885_in3)
          begin :bnn_N_Mux_2_4_8_1_1885
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1885_out1 = bnn_N_Mux_2_2_3_1_1807_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1885_out1 = bnn_N_Mux_2_4_8_1_1885_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1885_out1 = bnn_N_Mux_2_2_3_1_1810_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1885_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1885_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1886
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1886_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1886_out1 = bnn_N_Mux_2_4_8_1_1885_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1887_in3 = {bnn_RightShift_64Sx8S_1S_1_1728_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1886_out1 or bnn_N_Mux_2_2_3_1_1887_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1887
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1887_out1 = bnn_N_Mux_2_2_3_1_1886_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1887_out1 = bnn_N_Mux_2_2_3_1_1887_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1810_out1 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_N_Mux_2_4_8_1_1885_in3 or bnn_N_Mux_2_2_3_1_1887_out1)
          begin :bnn_N_Mux_2_4_8_1_1888
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1888_out1 = bnn_N_Mux_2_2_3_1_1887_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1888_out1 = bnn_N_Mux_2_4_8_1_1885_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1888_out1 = bnn_N_Mux_2_2_3_1_1810_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1888_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1888_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1889
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1889_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1889_out1 = bnn_N_Mux_2_4_8_1_1888_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1890_in3 = {bnn_RightShift_64Sx8S_1S_1_1648_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1889_out1 or bnn_N_Mux_2_2_3_1_1890_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1890
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1890_out1 = bnn_N_Mux_2_2_3_1_1889_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1890_out1 = bnn_N_Mux_2_2_3_1_1890_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1891_in1 = {s_reg_1076_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1891
         assign bnn_RightShift_64Sx8S_1S_1_1891_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1891_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1892_in3 = {bnn_RightShift_64Sx8S_1S_1_1891_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_937 or bnn_N_Mux_2_2_3_1_1892_in3)
          begin :bnn_N_Mux_2_2_3_1_1892
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1892_out1 = s_reg_937;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1892_out1 = bnn_N_Mux_2_2_3_1_1892_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_920 or s_reg_940 or s_reg_942 or bnn_N_Mux_2_2_3_1_1892_out1)
          begin :bnn_N_Mux_2_4_8_1_1893
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1893_out1 = bnn_N_Mux_2_2_3_1_1892_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1893_out1 = s_reg_940;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1893_out1 = s_reg_920;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1893_out1 = s_reg_942;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1893_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1894
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1894_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1894_out1 = bnn_N_Mux_2_4_8_1_1893_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1895_in3 = {bnn_RightShift_64Sx8S_1S_1_1705_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1894_out1 or bnn_N_Mux_2_2_3_1_1895_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1895
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1895_out1 = bnn_N_Mux_2_2_3_1_1894_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1895_out1 = bnn_N_Mux_2_2_3_1_1895_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1896_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[6], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1812_out1 or bnn_N_Mux_2_2_3_1_1815_out1 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_N_Mux_2_4_8_1_1896_in3)
          begin :bnn_N_Mux_2_4_8_1_1896
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1896_out1 = bnn_N_Mux_2_2_3_1_1812_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1896_out1 = bnn_N_Mux_2_4_8_1_1896_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1896_out1 = bnn_N_Mux_2_2_3_1_1815_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1896_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1896_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1897
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1897_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1897_out1 = bnn_N_Mux_2_4_8_1_1896_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1898_in3 = {bnn_RightShift_64Sx8S_1S_1_1729_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1897_out1 or bnn_N_Mux_2_2_3_1_1898_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1898
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1898_out1 = bnn_N_Mux_2_2_3_1_1897_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1898_out1 = bnn_N_Mux_2_2_3_1_1898_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1815_out1 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_N_Mux_2_4_8_1_1896_in3 or bnn_N_Mux_2_2_3_1_1898_out1)
          begin :bnn_N_Mux_2_4_8_1_1899
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1899_out1 = bnn_N_Mux_2_2_3_1_1898_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1899_out1 = bnn_N_Mux_2_4_8_1_1896_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1899_out1 = bnn_N_Mux_2_2_3_1_1815_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1899_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1899_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1900
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1900_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1900_out1 = bnn_N_Mux_2_4_8_1_1899_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1901_in3 = {bnn_RightShift_64Sx8S_1S_1_1649_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1900_out1 or bnn_N_Mux_2_2_3_1_1901_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1901
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1901_out1 = bnn_N_Mux_2_2_3_1_1900_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1901_out1 = bnn_N_Mux_2_2_3_1_1901_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1902_in1 = {s_reg_1076_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1902
         assign bnn_RightShift_64Sx8S_1S_1_1902_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1902_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1903_in3 = {bnn_RightShift_64Sx8S_1S_1_1902_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_941 or bnn_N_Mux_2_2_3_1_1903_in3)
          begin :bnn_N_Mux_2_2_3_1_1903
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1903_out1 = s_reg_941;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1903_out1 = bnn_N_Mux_2_2_3_1_1903_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_928 or s_reg_945 or s_reg_947 or bnn_N_Mux_2_2_3_1_1903_out1)
          begin :bnn_N_Mux_2_4_8_1_1904
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1904_out1 = bnn_N_Mux_2_2_3_1_1903_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1904_out1 = s_reg_945;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1904_out1 = s_reg_928;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1904_out1 = s_reg_947;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1904_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1905
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1905_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1905_out1 = bnn_N_Mux_2_4_8_1_1904_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1906_in3 = {bnn_RightShift_64Sx8S_1S_1_1706_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1905_out1 or bnn_N_Mux_2_2_3_1_1906_in3 or s_reg_1049_stage1)
          begin :bnn_N_Mux_2_2_3_1_1906
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1906_out1 = bnn_N_Mux_2_2_3_1_1905_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1906_out1 = bnn_N_Mux_2_2_3_1_1906_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1907_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[7], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1817_out1 or bnn_N_Mux_2_2_3_1_1820_out1 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_N_Mux_2_4_8_1_1907_in3)
          begin :bnn_N_Mux_2_4_8_1_1907
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1907_out1 = bnn_N_Mux_2_2_3_1_1817_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1907_out1 = bnn_N_Mux_2_4_8_1_1907_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1907_out1 = bnn_N_Mux_2_2_3_1_1820_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1907_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1907_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_1908
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_1908_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1908_out1 = bnn_N_Mux_2_4_8_1_1907_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1909_in3 = {bnn_RightShift_64Sx8S_1S_4_1730_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1908_out1 or bnn_N_Mux_2_2_3_1_1909_in3 or s_reg_1037_stage1)
          begin :bnn_N_Mux_2_2_3_1_1909
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_1909_out1 = bnn_N_Mux_2_2_3_1_1908_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1909_out1 = bnn_N_Mux_2_2_3_1_1909_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1820_out1 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_N_Mux_2_4_8_1_1907_in3 or bnn_N_Mux_2_2_3_1_1909_out1)
          begin :bnn_N_Mux_2_4_8_1_1910
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1910_out1 = bnn_N_Mux_2_2_3_1_1909_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1910_out1 = bnn_N_Mux_2_4_8_1_1907_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1910_out1 = bnn_N_Mux_2_2_3_1_1820_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1910_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1910_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_1911
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_1911_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1911_out1 = bnn_N_Mux_2_4_8_1_1910_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1912_in3 = {bnn_RightShift_64Sx8S_1S_4_1650_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1911_out1 or bnn_N_Mux_2_2_3_1_1912_in3 or s_reg_1038_stage1)
          begin :bnn_N_Mux_2_2_3_1_1912
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_1912_out1 = bnn_N_Mux_2_2_3_1_1911_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1912_out1 = bnn_N_Mux_2_2_3_1_1912_in3;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1913
         assign bnn_RightShift_64Sx8S_1S_1_1913_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1020_stage1_slice[5:0];

         assign bnn_N_Mux_3_2_6_1_1914_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_1913_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_1914_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_1914
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_1914_out1_slice = bnn_N_Mux_3_2_6_1_1914_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_1914_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_894 or bnn_N_Mux_3_2_6_1_1914_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1915
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_1915_out1 = s_reg_894;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1915_out1 = bnn_N_Mux_3_2_6_1_1914_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_891 or s_reg_902 or s_reg_905 or bnn_N_Mux_2_2_3_1_1915_out1)
          begin :bnn_N_Mux_2_4_8_1_1916
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1916_out1 = bnn_N_Mux_2_2_3_1_1915_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1916_out1 = s_reg_902;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1916_out1 = s_reg_891;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1916_out1 = s_reg_905;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1916_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_1917
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_1917_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1917_out1 = bnn_N_Mux_2_4_8_1_1916_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1917_out1 or s_reg_1049_stage1 or bnn_N_Mux_3_2_6_1_1698_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_1918
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_1918_out1 = bnn_N_Mux_2_2_3_1_1917_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1918_out1 = bnn_N_Mux_3_2_6_1_1698_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_7_4
         always @(s_reg_1004 or s_reg_879 or s_reg_883 or bnn_N_Mux_2_2_3_1_1918_out1)
          begin :bnn_N_Mux_2_4_7_4_1919
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_7_4_1919_out1 = s_reg_879;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_7_4_1919_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_7_4_1919_out1 = s_reg_883;
               end
               
               default: begin
                  bnn_N_Mux_2_4_7_4_1919_out1 = bnn_N_Mux_2_2_3_1_1918_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_1577_out1 or bnn_N_Mux_2_4_7_4_1919_out1)
          begin :bnn_N_Mux_3_2_6_4_1920
            if (bnn_And_1Sx1U_1U_4_1577_out1) begin
               bnn_N_Mux_3_2_6_4_1920_out1_slice = bnn_N_Mux_2_4_7_4_1919_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_1920_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_7_4
         always @(s_reg_1004 or s_reg_883 or bnn_N_Mux_2_2_3_1_1918_out1 or bnn_N_Mux_3_2_6_4_1920_out1_slice)
          begin :bnn_N_Mux_2_4_7_4_1921
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_7_4_1921_out1 = bnn_N_Mux_3_2_6_4_1920_out1_slice;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_7_4_1921_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_7_4_1921_out1 = s_reg_883;
               end
               
               default: begin
                  bnn_N_Mux_2_4_7_4_1921_out1 = bnn_N_Mux_2_2_3_1_1918_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_1578_out1 or bnn_N_Mux_2_4_7_4_1921_out1)
          begin :bnn_N_Mux_3_2_6_4_1922
            if (bnn_And_1Sx1U_1U_4_1578_out1) begin
               bnn_N_Mux_3_2_6_4_1922_out1_slice = bnn_N_Mux_2_4_7_4_1921_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_1922_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1923_in1 = {s_reg_1029_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1923
         assign bnn_RightShift_64Sx8S_1S_1_1923_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1923_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1924_in3 = {bnn_RightShift_64Sx8S_1S_1_1923_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_949 or bnn_N_Mux_2_2_3_1_1924_in3)
          begin :bnn_N_Mux_2_2_3_1_1924
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1924_out1 = s_reg_949;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1924_out1 = bnn_N_Mux_2_2_3_1_1924_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_896 or s_reg_954 or s_reg_956 or bnn_N_Mux_2_2_3_1_1924_out1)
          begin :bnn_N_Mux_2_4_8_1_1925
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1925_out1 = bnn_N_Mux_2_2_3_1_1924_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1925_out1 = s_reg_954;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1925_out1 = s_reg_896;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1925_out1 = s_reg_956;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1925_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1926
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1926_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1926_out1 = bnn_N_Mux_2_4_8_1_1925_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1927_in3 = {bnn_RightShift_64Sx8S_1S_1_1707_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1926_out1 or bnn_N_Mux_2_2_3_1_1927_in3)
          begin :bnn_N_Mux_2_2_3_1_1927
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1927_out1 = bnn_N_Mux_2_2_3_1_1926_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1927_out1 = bnn_N_Mux_2_2_3_1_1927_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1928_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[8], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1822_out1 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_N_Mux_2_4_8_1_1928_in3)
          begin :bnn_N_Mux_2_4_8_1_1928
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1928_out1 = bnn_N_Mux_2_2_3_1_1822_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1928_out1 = bnn_N_Mux_2_4_8_1_1928_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1928_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1928_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1928_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1929
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1929_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1929_out1 = bnn_N_Mux_2_4_8_1_1928_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1930_in3 = {bnn_RightShift_64Sx8S_1S_1_1731_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1929_out1 or bnn_N_Mux_2_2_3_1_1930_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1930
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1930_out1 = bnn_N_Mux_2_2_3_1_1929_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1930_out1 = bnn_N_Mux_2_2_3_1_1930_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_N_Mux_2_4_8_1_1928_in3 or bnn_N_Mux_2_2_3_1_1930_out1)
          begin :bnn_N_Mux_2_4_8_1_1931
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1931_out1 = bnn_N_Mux_2_2_3_1_1930_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1931_out1 = bnn_N_Mux_2_4_8_1_1928_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1931_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1931_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1931_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1932
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1932_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1932_out1 = bnn_N_Mux_2_4_8_1_1931_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1933_in3 = {bnn_RightShift_64Sx8S_1S_1_1651_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1932_out1 or bnn_N_Mux_2_2_3_1_1933_in3)
          begin :bnn_N_Mux_2_2_3_1_1933
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1933_out1 = bnn_N_Mux_2_2_3_1_1932_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1933_out1 = bnn_N_Mux_2_2_3_1_1933_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1934_in1 = {s_reg_1029_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1934
         assign bnn_RightShift_64Sx8S_1S_1_1934_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1934_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1935_in3 = {bnn_RightShift_64Sx8S_1S_1_1934_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_955 or bnn_N_Mux_2_2_3_1_1935_in3)
          begin :bnn_N_Mux_2_2_3_1_1935
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1935_out1 = s_reg_955;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1935_out1 = bnn_N_Mux_2_2_3_1_1935_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_906 or s_reg_958 or s_reg_960 or bnn_N_Mux_2_2_3_1_1935_out1)
          begin :bnn_N_Mux_2_4_8_1_1936
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1936_out1 = bnn_N_Mux_2_2_3_1_1935_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1936_out1 = s_reg_958;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1936_out1 = s_reg_906;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1936_out1 = s_reg_960;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1936_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1937
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1937_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1937_out1 = bnn_N_Mux_2_4_8_1_1936_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1938_in3 = {bnn_RightShift_64Sx8S_1S_1_1708_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1937_out1 or bnn_N_Mux_2_2_3_1_1938_in3)
          begin :bnn_N_Mux_2_2_3_1_1938
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1938_out1 = bnn_N_Mux_2_2_3_1_1937_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1938_out1 = bnn_N_Mux_2_2_3_1_1938_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1939_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[9], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1837_out1 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_N_Mux_2_4_8_1_1939_in3)
          begin :bnn_N_Mux_2_4_8_1_1939
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1939_out1 = bnn_N_Mux_2_2_3_1_1837_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1939_out1 = bnn_N_Mux_2_4_8_1_1939_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1939_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1939_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1939_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1940
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1940_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1940_out1 = bnn_N_Mux_2_4_8_1_1939_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1941_in3 = {bnn_RightShift_64Sx8S_1S_1_1732_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1940_out1 or bnn_N_Mux_2_2_3_1_1941_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1941
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1941_out1 = bnn_N_Mux_2_2_3_1_1940_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1941_out1 = bnn_N_Mux_2_2_3_1_1941_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_N_Mux_2_4_8_1_1939_in3 or bnn_N_Mux_2_2_3_1_1941_out1)
          begin :bnn_N_Mux_2_4_8_1_1942
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1942_out1 = bnn_N_Mux_2_2_3_1_1941_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1942_out1 = bnn_N_Mux_2_4_8_1_1939_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1942_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1942_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1942_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1943
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1943_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1943_out1 = bnn_N_Mux_2_4_8_1_1942_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1944_in3 = {bnn_RightShift_64Sx8S_1S_1_1652_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1943_out1 or bnn_N_Mux_2_2_3_1_1944_in3)
          begin :bnn_N_Mux_2_2_3_1_1944
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1944_out1 = bnn_N_Mux_2_2_3_1_1943_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1944_out1 = bnn_N_Mux_2_2_3_1_1944_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1945_in1 = {s_reg_1029_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1945
         assign bnn_RightShift_64Sx8S_1S_1_1945_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1945_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1946_in3 = {bnn_RightShift_64Sx8S_1S_1_1945_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_959 or bnn_N_Mux_2_2_3_1_1946_in3)
          begin :bnn_N_Mux_2_2_3_1_1946
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1946_out1 = s_reg_959;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1946_out1 = bnn_N_Mux_2_2_3_1_1946_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_915 or s_reg_961 or s_reg_963 or bnn_N_Mux_2_2_3_1_1946_out1)
          begin :bnn_N_Mux_2_4_8_1_1947
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1947_out1 = bnn_N_Mux_2_2_3_1_1946_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1947_out1 = s_reg_961;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1947_out1 = s_reg_915;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1947_out1 = s_reg_963;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1947_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1948
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1948_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1948_out1 = bnn_N_Mux_2_4_8_1_1947_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1949_in3 = {bnn_RightShift_64Sx8S_1S_1_1709_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1948_out1 or bnn_N_Mux_2_2_3_1_1949_in3)
          begin :bnn_N_Mux_2_2_3_1_1949
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1949_out1 = bnn_N_Mux_2_2_3_1_1948_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1949_out1 = bnn_N_Mux_2_2_3_1_1949_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1950_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[10], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1848_out1 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_N_Mux_2_4_8_1_1950_in3)
          begin :bnn_N_Mux_2_4_8_1_1950
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1950_out1 = bnn_N_Mux_2_2_3_1_1848_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1950_out1 = bnn_N_Mux_2_4_8_1_1950_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1950_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1950_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1950_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1951
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1951_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1951_out1 = bnn_N_Mux_2_4_8_1_1950_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1952_in3 = {bnn_RightShift_64Sx8S_1S_1_1733_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1951_out1 or bnn_N_Mux_2_2_3_1_1952_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1952
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1952_out1 = bnn_N_Mux_2_2_3_1_1951_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1952_out1 = bnn_N_Mux_2_2_3_1_1952_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_N_Mux_2_4_8_1_1950_in3 or bnn_N_Mux_2_2_3_1_1952_out1)
          begin :bnn_N_Mux_2_4_8_1_1953
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1953_out1 = bnn_N_Mux_2_2_3_1_1952_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1953_out1 = bnn_N_Mux_2_4_8_1_1950_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1953_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1953_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1953_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1954
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1954_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1954_out1 = bnn_N_Mux_2_4_8_1_1953_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1955_in3 = {bnn_RightShift_64Sx8S_1S_1_1653_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1954_out1 or bnn_N_Mux_2_2_3_1_1955_in3)
          begin :bnn_N_Mux_2_2_3_1_1955
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1955_out1 = bnn_N_Mux_2_2_3_1_1954_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1955_out1 = bnn_N_Mux_2_2_3_1_1955_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1956_in1 = {s_reg_1029_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1956
         assign bnn_RightShift_64Sx8S_1S_1_1956_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1956_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1957_in3 = {bnn_RightShift_64Sx8S_1S_1_1956_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_962 or bnn_N_Mux_2_2_3_1_1957_in3)
          begin :bnn_N_Mux_2_2_3_1_1957
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1957_out1 = s_reg_962;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1957_out1 = bnn_N_Mux_2_2_3_1_1957_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_923 or s_reg_964 or s_reg_966 or bnn_N_Mux_2_2_3_1_1957_out1)
          begin :bnn_N_Mux_2_4_8_1_1958
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1958_out1 = bnn_N_Mux_2_2_3_1_1957_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1958_out1 = s_reg_964;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1958_out1 = s_reg_923;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1958_out1 = s_reg_966;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1958_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1959
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1959_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1959_out1 = bnn_N_Mux_2_4_8_1_1958_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1960_in3 = {bnn_RightShift_64Sx8S_1S_1_1710_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1959_out1 or bnn_N_Mux_2_2_3_1_1960_in3)
          begin :bnn_N_Mux_2_2_3_1_1960
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1960_out1 = bnn_N_Mux_2_2_3_1_1959_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1960_out1 = bnn_N_Mux_2_2_3_1_1960_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1961_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[11], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1859_out1 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_N_Mux_2_4_8_1_1961_in3)
          begin :bnn_N_Mux_2_4_8_1_1961
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1961_out1 = bnn_N_Mux_2_2_3_1_1859_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1961_out1 = bnn_N_Mux_2_4_8_1_1961_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1961_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1961_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1961_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1962
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1962_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1962_out1 = bnn_N_Mux_2_4_8_1_1961_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1963_in3 = {bnn_RightShift_64Sx8S_1S_1_1734_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1962_out1 or bnn_N_Mux_2_2_3_1_1963_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1963
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1963_out1 = bnn_N_Mux_2_2_3_1_1962_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1963_out1 = bnn_N_Mux_2_2_3_1_1963_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_N_Mux_2_4_8_1_1961_in3 or bnn_N_Mux_2_2_3_1_1963_out1)
          begin :bnn_N_Mux_2_4_8_1_1964
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1964_out1 = bnn_N_Mux_2_2_3_1_1963_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1964_out1 = bnn_N_Mux_2_4_8_1_1961_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1964_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1964_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1964_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1965
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1965_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1965_out1 = bnn_N_Mux_2_4_8_1_1964_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1966_in3 = {bnn_RightShift_64Sx8S_1S_1_1654_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1965_out1 or bnn_N_Mux_2_2_3_1_1966_in3)
          begin :bnn_N_Mux_2_2_3_1_1966
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1966_out1 = bnn_N_Mux_2_2_3_1_1965_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1966_out1 = bnn_N_Mux_2_2_3_1_1966_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1967_in1 = {s_reg_1029_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1967
         assign bnn_RightShift_64Sx8S_1S_1_1967_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1967_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1968_in3 = {bnn_RightShift_64Sx8S_1S_1_1967_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_965 or bnn_N_Mux_2_2_3_1_1968_in3)
          begin :bnn_N_Mux_2_2_3_1_1968
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1968_out1 = s_reg_965;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1968_out1 = bnn_N_Mux_2_2_3_1_1968_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_931 or s_reg_967 or s_reg_969 or bnn_N_Mux_2_2_3_1_1968_out1)
          begin :bnn_N_Mux_2_4_8_1_1969
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1969_out1 = bnn_N_Mux_2_2_3_1_1968_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1969_out1 = s_reg_967;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1969_out1 = s_reg_931;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1969_out1 = s_reg_969;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1969_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1970
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1970_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1970_out1 = bnn_N_Mux_2_4_8_1_1969_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1971_in3 = {bnn_RightShift_64Sx8S_1S_1_1711_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1970_out1 or bnn_N_Mux_2_2_3_1_1971_in3)
          begin :bnn_N_Mux_2_2_3_1_1971
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1971_out1 = bnn_N_Mux_2_2_3_1_1970_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1971_out1 = bnn_N_Mux_2_2_3_1_1971_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1972_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[12], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1870_out1 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_N_Mux_2_4_8_1_1972_in3)
          begin :bnn_N_Mux_2_4_8_1_1972
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1972_out1 = bnn_N_Mux_2_2_3_1_1870_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1972_out1 = bnn_N_Mux_2_4_8_1_1972_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1972_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1972_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1972_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1973
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1973_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1973_out1 = bnn_N_Mux_2_4_8_1_1972_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1974_in3 = {bnn_RightShift_64Sx8S_1S_1_1735_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1973_out1 or bnn_N_Mux_2_2_3_1_1974_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1974
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1974_out1 = bnn_N_Mux_2_2_3_1_1973_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1974_out1 = bnn_N_Mux_2_2_3_1_1974_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_N_Mux_2_4_8_1_1972_in3 or bnn_N_Mux_2_2_3_1_1974_out1)
          begin :bnn_N_Mux_2_4_8_1_1975
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1975_out1 = bnn_N_Mux_2_2_3_1_1974_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1975_out1 = bnn_N_Mux_2_4_8_1_1972_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1975_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1975_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1975_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1976
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1976_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1976_out1 = bnn_N_Mux_2_4_8_1_1975_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1977_in3 = {bnn_RightShift_64Sx8S_1S_1_1655_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1976_out1 or bnn_N_Mux_2_2_3_1_1977_in3)
          begin :bnn_N_Mux_2_2_3_1_1977
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1977_out1 = bnn_N_Mux_2_2_3_1_1976_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1977_out1 = bnn_N_Mux_2_2_3_1_1977_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1978_in1 = {s_reg_1029_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1978
         assign bnn_RightShift_64Sx8S_1S_1_1978_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1978_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1979_in3 = {bnn_RightShift_64Sx8S_1S_1_1978_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_968 or bnn_N_Mux_2_2_3_1_1979_in3)
          begin :bnn_N_Mux_2_2_3_1_1979
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1979_out1 = s_reg_968;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1979_out1 = bnn_N_Mux_2_2_3_1_1979_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_938 or s_reg_970 or s_reg_972 or bnn_N_Mux_2_2_3_1_1979_out1)
          begin :bnn_N_Mux_2_4_8_1_1980
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1980_out1 = bnn_N_Mux_2_2_3_1_1979_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1980_out1 = s_reg_970;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1980_out1 = s_reg_938;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1980_out1 = s_reg_972;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1980_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1981
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1981_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1981_out1 = bnn_N_Mux_2_4_8_1_1980_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1982_in3 = {bnn_RightShift_64Sx8S_1S_1_1712_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1981_out1 or bnn_N_Mux_2_2_3_1_1982_in3)
          begin :bnn_N_Mux_2_2_3_1_1982
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1982_out1 = bnn_N_Mux_2_2_3_1_1981_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1982_out1 = bnn_N_Mux_2_2_3_1_1982_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1983_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[13], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1881_out1 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_N_Mux_2_4_8_1_1983_in3)
          begin :bnn_N_Mux_2_4_8_1_1983
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1983_out1 = bnn_N_Mux_2_2_3_1_1881_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1983_out1 = bnn_N_Mux_2_4_8_1_1983_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1983_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1983_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1983_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1984
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1984_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1984_out1 = bnn_N_Mux_2_4_8_1_1983_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1985_in3 = {bnn_RightShift_64Sx8S_1S_1_1736_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1984_out1 or bnn_N_Mux_2_2_3_1_1985_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1985
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1985_out1 = bnn_N_Mux_2_2_3_1_1984_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1985_out1 = bnn_N_Mux_2_2_3_1_1985_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_N_Mux_2_4_8_1_1983_in3 or bnn_N_Mux_2_2_3_1_1985_out1)
          begin :bnn_N_Mux_2_4_8_1_1986
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1986_out1 = bnn_N_Mux_2_2_3_1_1985_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1986_out1 = bnn_N_Mux_2_4_8_1_1983_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1986_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1986_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1986_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1987
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1987_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1987_out1 = bnn_N_Mux_2_4_8_1_1986_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1988_in3 = {bnn_RightShift_64Sx8S_1S_1_1656_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1987_out1 or bnn_N_Mux_2_2_3_1_1988_in3)
          begin :bnn_N_Mux_2_2_3_1_1988
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1988_out1 = bnn_N_Mux_2_2_3_1_1987_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1988_out1 = bnn_N_Mux_2_2_3_1_1988_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_1989_in1 = {s_reg_1029_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_1989
         assign bnn_RightShift_64Sx8S_1S_1_1989_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_1989_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_1990_in3 = {bnn_RightShift_64Sx8S_1S_1_1989_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_971 or bnn_N_Mux_2_2_3_1_1990_in3)
          begin :bnn_N_Mux_2_2_3_1_1990
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_1990_out1 = s_reg_971;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1990_out1 = bnn_N_Mux_2_2_3_1_1990_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_942 or s_reg_973 or s_reg_975 or bnn_N_Mux_2_2_3_1_1990_out1)
          begin :bnn_N_Mux_2_4_8_1_1991
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1991_out1 = bnn_N_Mux_2_2_3_1_1990_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1991_out1 = s_reg_973;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1991_out1 = s_reg_942;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1991_out1 = s_reg_975;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1991_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_1992
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_1992_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1992_out1 = bnn_N_Mux_2_4_8_1_1991_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1993_in3 = {bnn_RightShift_64Sx8S_1S_1_1713_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_1992_out1 or bnn_N_Mux_2_2_3_1_1993_in3)
          begin :bnn_N_Mux_2_2_3_1_1993
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_1993_out1 = bnn_N_Mux_2_2_3_1_1992_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1993_out1 = bnn_N_Mux_2_2_3_1_1993_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_1994_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[14], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1892_out1 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_N_Mux_2_4_8_1_1994_in3)
          begin :bnn_N_Mux_2_4_8_1_1994
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1994_out1 = bnn_N_Mux_2_2_3_1_1892_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1994_out1 = bnn_N_Mux_2_4_8_1_1994_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1994_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1994_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1994_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_1995
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_1995_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1995_out1 = bnn_N_Mux_2_4_8_1_1994_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1996_in3 = {bnn_RightShift_64Sx8S_1S_1_1737_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_1995_out1 or bnn_N_Mux_2_2_3_1_1996_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_1996
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_1996_out1 = bnn_N_Mux_2_2_3_1_1995_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1996_out1 = bnn_N_Mux_2_2_3_1_1996_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_N_Mux_2_4_8_1_1994_in3 or bnn_N_Mux_2_2_3_1_1996_out1)
          begin :bnn_N_Mux_2_4_8_1_1997
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_1997_out1 = bnn_N_Mux_2_2_3_1_1996_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_1997_out1 = bnn_N_Mux_2_4_8_1_1994_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_1997_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_1997_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_1997_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_1998
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_1998_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1998_out1 = bnn_N_Mux_2_4_8_1_1997_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_1999_in3 = {bnn_RightShift_64Sx8S_1S_1_1657_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_1998_out1 or bnn_N_Mux_2_2_3_1_1999_in3)
          begin :bnn_N_Mux_2_2_3_1_1999
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_1999_out1 = bnn_N_Mux_2_2_3_1_1998_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_1999_out1 = bnn_N_Mux_2_2_3_1_1999_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2000_in1 = {s_reg_1029_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2000
         assign bnn_RightShift_64Sx8S_1S_1_2000_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2000_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2001_in3 = {bnn_RightShift_64Sx8S_1S_1_2000_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_974 or bnn_N_Mux_2_2_3_1_2001_in3)
          begin :bnn_N_Mux_2_2_3_1_2001
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_2001_out1 = s_reg_974;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2001_out1 = bnn_N_Mux_2_2_3_1_2001_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_947 or s_reg_978 or s_reg_980 or bnn_N_Mux_2_2_3_1_2001_out1)
          begin :bnn_N_Mux_2_4_8_1_2002
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2002_out1 = bnn_N_Mux_2_2_3_1_2001_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2002_out1 = s_reg_978;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2002_out1 = s_reg_947;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2002_out1 = s_reg_980;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2002_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_2003
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_2003_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2003_out1 = bnn_N_Mux_2_4_8_1_2002_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2004_in3 = {bnn_RightShift_64Sx8S_1S_1_1714_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_2003_out1 or bnn_N_Mux_2_2_3_1_2004_in3)
          begin :bnn_N_Mux_2_2_3_1_2004
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_2004_out1 = bnn_N_Mux_2_2_3_1_2003_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2004_out1 = bnn_N_Mux_2_2_3_1_2004_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2005_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[15], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1903_out1 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_N_Mux_2_4_8_1_2005_in3)
          begin :bnn_N_Mux_2_4_8_1_2005
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2005_out1 = bnn_N_Mux_2_2_3_1_1903_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2005_out1 = bnn_N_Mux_2_4_8_1_2005_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2005_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2005_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2005_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_2006
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_2006_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2006_out1 = bnn_N_Mux_2_4_8_1_2005_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2007_in3 = {bnn_RightShift_64Sx8S_1S_1_1738_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2006_out1 or bnn_N_Mux_2_2_3_1_2007_in3 or s_reg_1051_stage1)
          begin :bnn_N_Mux_2_2_3_1_2007
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_2007_out1 = bnn_N_Mux_2_2_3_1_2006_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2007_out1 = bnn_N_Mux_2_2_3_1_2007_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_N_Mux_2_4_8_1_2005_in3 or bnn_N_Mux_2_2_3_1_2007_out1)
          begin :bnn_N_Mux_2_4_8_1_2008
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2008_out1 = bnn_N_Mux_2_2_3_1_2007_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2008_out1 = bnn_N_Mux_2_4_8_1_2005_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2008_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2008_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2008_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_2009
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_2009_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2009_out1 = bnn_N_Mux_2_4_8_1_2008_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2010_in3 = {bnn_RightShift_64Sx8S_1S_1_1658_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_2009_out1 or bnn_N_Mux_2_2_3_1_2010_in3)
          begin :bnn_N_Mux_2_2_3_1_2010
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_2010_out1 = bnn_N_Mux_2_2_3_1_2009_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2010_out1 = bnn_N_Mux_2_2_3_1_2010_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2011_in1 = {s_reg_1093_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2011
         assign bnn_RightShift_64Sx8S_1S_1_2011_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2011_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2012_in3 = {bnn_RightShift_64Sx8S_1S_1_2011_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_982 or bnn_N_Mux_2_2_3_1_2012_in3)
          begin :bnn_N_Mux_2_2_3_1_2012
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2012_out1 = s_reg_982;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2012_out1 = bnn_N_Mux_2_2_3_1_2012_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_956 or s_reg_977 or s_reg_985 or bnn_N_Mux_2_2_3_1_2012_out1)
          begin :bnn_N_Mux_2_4_8_1_2013
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2013_out1 = bnn_N_Mux_2_2_3_1_2012_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2013_out1 = s_reg_985;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2013_out1 = s_reg_956;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2013_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2013_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2014
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2014_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2014_out1 = bnn_N_Mux_2_4_8_1_2013_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2015_in3 = {bnn_RightShift_64Sx8S_1S_1_1715_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2014_out1 or bnn_N_Mux_2_2_3_1_2015_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2015
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2015_out1 = bnn_N_Mux_2_2_3_1_2014_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2015_out1 = bnn_N_Mux_2_2_3_1_2015_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2016_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[16], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1924_out1 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_N_Mux_2_4_8_1_2016_in3)
          begin :bnn_N_Mux_2_4_8_1_2016
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2016_out1 = bnn_N_Mux_2_2_3_1_1924_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2016_out1 = bnn_N_Mux_2_4_8_1_2016_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2016_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2016_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2016_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2017
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2017_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2017_out1 = bnn_N_Mux_2_4_8_1_2016_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2018_in3 = {bnn_RightShift_64Sx8S_1S_1_1739_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2017_out1 or bnn_N_Mux_2_2_3_1_2018_in3)
          begin :bnn_N_Mux_2_2_3_1_2018
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2018_out1 = bnn_N_Mux_2_2_3_1_2017_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2018_out1 = bnn_N_Mux_2_2_3_1_2018_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_N_Mux_2_4_8_1_2016_in3 or bnn_N_Mux_2_2_3_1_2018_out1)
          begin :bnn_N_Mux_2_4_8_1_2019
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2019_out1 = bnn_N_Mux_2_2_3_1_2018_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2019_out1 = bnn_N_Mux_2_4_8_1_2016_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2019_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2019_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2019_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2020
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2020_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2020_out1 = bnn_N_Mux_2_4_8_1_2019_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2021_in3 = {bnn_RightShift_64Sx8S_1S_1_1659_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2020_out1 or bnn_N_Mux_2_2_3_1_2021_in3)
          begin :bnn_N_Mux_2_2_3_1_2021
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2021_out1 = bnn_N_Mux_2_2_3_1_2020_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2021_out1 = bnn_N_Mux_2_2_3_1_2021_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2022_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[24], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2012_out1 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_N_Mux_2_4_8_1_2022_in3)
          begin :bnn_N_Mux_2_4_8_1_2022
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2022_out1 = bnn_N_Mux_2_2_3_1_2012_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2022_out1 = bnn_N_Mux_2_4_8_1_2022_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2022_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2022_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2022_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2023
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2023_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2023_out1 = bnn_N_Mux_2_4_8_1_2022_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2024_in3 = {bnn_RightShift_64Sx8S_1S_1_1747_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2023_out1 or bnn_N_Mux_2_2_3_1_2024_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2024
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2024_out1 = bnn_N_Mux_2_2_3_1_2023_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2024_out1 = bnn_N_Mux_2_2_3_1_2024_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_N_Mux_2_4_8_1_2022_in3 or bnn_N_Mux_2_2_3_1_2024_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2025
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2025_out1 = bnn_N_Mux_2_2_3_1_2024_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2025_out1 = bnn_N_Mux_2_4_8_1_2022_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2025_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2025_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2025_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2026
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2026_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2026_out1 = bnn_N_Mux_2_4_8_1_2025_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2027_in3 = {bnn_RightShift_64Sx8S_1S_1_1667_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2026_out1 or bnn_N_Mux_2_2_3_1_2027_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2027
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2027_out1 = bnn_N_Mux_2_2_3_1_2026_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2027_out1 = bnn_N_Mux_2_2_3_1_2027_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2028_in1 = {s_reg_1093_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2028
         assign bnn_RightShift_64Sx8S_1S_1_2028_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2028_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2029_in3 = {bnn_RightShift_64Sx8S_1S_1_2028_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_986 or bnn_N_Mux_2_2_3_1_2029_in3)
          begin :bnn_N_Mux_2_2_3_1_2029
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2029_out1 = s_reg_986;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2029_out1 = bnn_N_Mux_2_2_3_1_2029_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_960 or s_reg_977 or s_reg_987 or bnn_N_Mux_2_2_3_1_2029_out1)
          begin :bnn_N_Mux_2_4_8_1_2030
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2030_out1 = bnn_N_Mux_2_2_3_1_2029_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2030_out1 = s_reg_987;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2030_out1 = s_reg_960;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2030_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2030_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2031
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2031_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2031_out1 = bnn_N_Mux_2_4_8_1_2030_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2032_in3 = {bnn_RightShift_64Sx8S_1S_1_1716_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2031_out1 or bnn_N_Mux_2_2_3_1_2032_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2032
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2032_out1 = bnn_N_Mux_2_2_3_1_2031_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2032_out1 = bnn_N_Mux_2_2_3_1_2032_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2033_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[17], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1935_out1 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_N_Mux_2_4_8_1_2033_in3)
          begin :bnn_N_Mux_2_4_8_1_2033
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2033_out1 = bnn_N_Mux_2_2_3_1_1935_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2033_out1 = bnn_N_Mux_2_4_8_1_2033_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2033_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2033_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2033_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2034
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2034_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2034_out1 = bnn_N_Mux_2_4_8_1_2033_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2035_in3 = {bnn_RightShift_64Sx8S_1S_1_1740_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2034_out1 or bnn_N_Mux_2_2_3_1_2035_in3)
          begin :bnn_N_Mux_2_2_3_1_2035
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2035_out1 = bnn_N_Mux_2_2_3_1_2034_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2035_out1 = bnn_N_Mux_2_2_3_1_2035_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_N_Mux_2_4_8_1_2033_in3 or bnn_N_Mux_2_2_3_1_2035_out1)
          begin :bnn_N_Mux_2_4_8_1_2036
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2036_out1 = bnn_N_Mux_2_2_3_1_2035_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2036_out1 = bnn_N_Mux_2_4_8_1_2033_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2036_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2036_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2036_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2037
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2037_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2037_out1 = bnn_N_Mux_2_4_8_1_2036_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2038_in3 = {bnn_RightShift_64Sx8S_1S_1_1660_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2037_out1 or bnn_N_Mux_2_2_3_1_2038_in3)
          begin :bnn_N_Mux_2_2_3_1_2038
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2038_out1 = bnn_N_Mux_2_2_3_1_2037_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2038_out1 = bnn_N_Mux_2_2_3_1_2038_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2039_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[25], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2029_out1 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_N_Mux_2_4_8_1_2039_in3)
          begin :bnn_N_Mux_2_4_8_1_2039
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2039_out1 = bnn_N_Mux_2_2_3_1_2029_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2039_out1 = bnn_N_Mux_2_4_8_1_2039_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2039_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2039_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2039_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2040
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2040_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2040_out1 = bnn_N_Mux_2_4_8_1_2039_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2041_in3 = {bnn_RightShift_64Sx8S_1S_1_1748_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2040_out1 or bnn_N_Mux_2_2_3_1_2041_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2041
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2041_out1 = bnn_N_Mux_2_2_3_1_2040_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2041_out1 = bnn_N_Mux_2_2_3_1_2041_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_N_Mux_2_4_8_1_2039_in3 or bnn_N_Mux_2_2_3_1_2041_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2042
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2042_out1 = bnn_N_Mux_2_2_3_1_2041_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2042_out1 = bnn_N_Mux_2_4_8_1_2039_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2042_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2042_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2042_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2043
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2043_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2043_out1 = bnn_N_Mux_2_4_8_1_2042_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2044_in3 = {bnn_RightShift_64Sx8S_1S_1_1668_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2043_out1 or bnn_N_Mux_2_2_3_1_2044_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2044
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2044_out1 = bnn_N_Mux_2_2_3_1_2043_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2044_out1 = bnn_N_Mux_2_2_3_1_2044_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2045_in1 = {s_reg_1093_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2045
         assign bnn_RightShift_64Sx8S_1S_1_2045_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2045_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2046_in3 = {bnn_RightShift_64Sx8S_1S_1_2045_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_988 or bnn_N_Mux_2_2_3_1_2046_in3)
          begin :bnn_N_Mux_2_2_3_1_2046
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2046_out1 = s_reg_988;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2046_out1 = bnn_N_Mux_2_2_3_1_2046_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_963 or s_reg_977 or s_reg_989 or bnn_N_Mux_2_2_3_1_2046_out1)
          begin :bnn_N_Mux_2_4_8_1_2047
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2047_out1 = bnn_N_Mux_2_2_3_1_2046_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2047_out1 = s_reg_989;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2047_out1 = s_reg_963;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2047_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2047_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2048
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2048_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2048_out1 = bnn_N_Mux_2_4_8_1_2047_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2049_in3 = {bnn_RightShift_64Sx8S_1S_1_1717_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2048_out1 or bnn_N_Mux_2_2_3_1_2049_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2049
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2049_out1 = bnn_N_Mux_2_2_3_1_2048_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2049_out1 = bnn_N_Mux_2_2_3_1_2049_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2050_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[18], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1946_out1 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_N_Mux_2_4_8_1_2050_in3)
          begin :bnn_N_Mux_2_4_8_1_2050
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2050_out1 = bnn_N_Mux_2_2_3_1_1946_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2050_out1 = bnn_N_Mux_2_4_8_1_2050_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2050_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2050_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2050_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2051
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2051_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2051_out1 = bnn_N_Mux_2_4_8_1_2050_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2052_in3 = {bnn_RightShift_64Sx8S_1S_1_1741_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2051_out1 or bnn_N_Mux_2_2_3_1_2052_in3)
          begin :bnn_N_Mux_2_2_3_1_2052
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2052_out1 = bnn_N_Mux_2_2_3_1_2051_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2052_out1 = bnn_N_Mux_2_2_3_1_2052_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_N_Mux_2_4_8_1_2050_in3 or bnn_N_Mux_2_2_3_1_2052_out1)
          begin :bnn_N_Mux_2_4_8_1_2053
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2053_out1 = bnn_N_Mux_2_2_3_1_2052_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2053_out1 = bnn_N_Mux_2_4_8_1_2050_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2053_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2053_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2053_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2054
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2054_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2054_out1 = bnn_N_Mux_2_4_8_1_2053_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2055_in3 = {bnn_RightShift_64Sx8S_1S_1_1661_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2054_out1 or bnn_N_Mux_2_2_3_1_2055_in3)
          begin :bnn_N_Mux_2_2_3_1_2055
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2055_out1 = bnn_N_Mux_2_2_3_1_2054_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2055_out1 = bnn_N_Mux_2_2_3_1_2055_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2056_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[26], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2046_out1 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_N_Mux_2_4_8_1_2056_in3)
          begin :bnn_N_Mux_2_4_8_1_2056
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2056_out1 = bnn_N_Mux_2_2_3_1_2046_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2056_out1 = bnn_N_Mux_2_4_8_1_2056_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2056_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2056_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2056_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2057
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2057_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2057_out1 = bnn_N_Mux_2_4_8_1_2056_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2058_in3 = {bnn_RightShift_64Sx8S_1S_1_1749_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2057_out1 or bnn_N_Mux_2_2_3_1_2058_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2058
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2058_out1 = bnn_N_Mux_2_2_3_1_2057_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2058_out1 = bnn_N_Mux_2_2_3_1_2058_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_N_Mux_2_4_8_1_2056_in3 or bnn_N_Mux_2_2_3_1_2058_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2059
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2059_out1 = bnn_N_Mux_2_2_3_1_2058_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2059_out1 = bnn_N_Mux_2_4_8_1_2056_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2059_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2059_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2059_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2060
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2060_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2060_out1 = bnn_N_Mux_2_4_8_1_2059_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2061_in3 = {bnn_RightShift_64Sx8S_1S_1_1669_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2060_out1 or bnn_N_Mux_2_2_3_1_2061_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2061
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2061_out1 = bnn_N_Mux_2_2_3_1_2060_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2061_out1 = bnn_N_Mux_2_2_3_1_2061_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2062_in1 = {s_reg_1093_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2062
         assign bnn_RightShift_64Sx8S_1S_1_2062_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2062_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2063_in3 = {bnn_RightShift_64Sx8S_1S_1_2062_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_990 or bnn_N_Mux_2_2_3_1_2063_in3)
          begin :bnn_N_Mux_2_2_3_1_2063
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2063_out1 = s_reg_990;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2063_out1 = bnn_N_Mux_2_2_3_1_2063_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_966 or s_reg_977 or s_reg_991 or bnn_N_Mux_2_2_3_1_2063_out1)
          begin :bnn_N_Mux_2_4_8_1_2064
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2064_out1 = bnn_N_Mux_2_2_3_1_2063_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2064_out1 = s_reg_991;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2064_out1 = s_reg_966;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2064_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2064_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2065
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2065_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2065_out1 = bnn_N_Mux_2_4_8_1_2064_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2066_in3 = {bnn_RightShift_64Sx8S_1S_1_1718_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2065_out1 or bnn_N_Mux_2_2_3_1_2066_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2066
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2066_out1 = bnn_N_Mux_2_2_3_1_2065_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2066_out1 = bnn_N_Mux_2_2_3_1_2066_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2067_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[19], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1957_out1 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_N_Mux_2_4_8_1_2067_in3)
          begin :bnn_N_Mux_2_4_8_1_2067
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2067_out1 = bnn_N_Mux_2_2_3_1_1957_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2067_out1 = bnn_N_Mux_2_4_8_1_2067_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2067_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2067_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2067_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2068
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2068_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2068_out1 = bnn_N_Mux_2_4_8_1_2067_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2069_in3 = {bnn_RightShift_64Sx8S_1S_1_1742_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2068_out1 or bnn_N_Mux_2_2_3_1_2069_in3)
          begin :bnn_N_Mux_2_2_3_1_2069
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2069_out1 = bnn_N_Mux_2_2_3_1_2068_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2069_out1 = bnn_N_Mux_2_2_3_1_2069_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_N_Mux_2_4_8_1_2067_in3 or bnn_N_Mux_2_2_3_1_2069_out1)
          begin :bnn_N_Mux_2_4_8_1_2070
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2070_out1 = bnn_N_Mux_2_2_3_1_2069_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2070_out1 = bnn_N_Mux_2_4_8_1_2067_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2070_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2070_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2070_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2071
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2071_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2071_out1 = bnn_N_Mux_2_4_8_1_2070_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2072_in3 = {bnn_RightShift_64Sx8S_1S_1_1662_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2071_out1 or bnn_N_Mux_2_2_3_1_2072_in3)
          begin :bnn_N_Mux_2_2_3_1_2072
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2072_out1 = bnn_N_Mux_2_2_3_1_2071_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2072_out1 = bnn_N_Mux_2_2_3_1_2072_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2073_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[27], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2063_out1 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_N_Mux_2_4_8_1_2073_in3)
          begin :bnn_N_Mux_2_4_8_1_2073
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2073_out1 = bnn_N_Mux_2_2_3_1_2063_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2073_out1 = bnn_N_Mux_2_4_8_1_2073_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2073_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2073_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2073_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2074
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2074_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2074_out1 = bnn_N_Mux_2_4_8_1_2073_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2075_in3 = {bnn_RightShift_64Sx8S_1S_1_1750_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2074_out1 or bnn_N_Mux_2_2_3_1_2075_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2075
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2075_out1 = bnn_N_Mux_2_2_3_1_2074_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2075_out1 = bnn_N_Mux_2_2_3_1_2075_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_N_Mux_2_4_8_1_2073_in3 or bnn_N_Mux_2_2_3_1_2075_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2076
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2076_out1 = bnn_N_Mux_2_2_3_1_2075_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2076_out1 = bnn_N_Mux_2_4_8_1_2073_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2076_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2076_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2076_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2077
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2077_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2077_out1 = bnn_N_Mux_2_4_8_1_2076_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2078_in3 = {bnn_RightShift_64Sx8S_1S_1_1670_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2077_out1 or bnn_N_Mux_2_2_3_1_2078_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2078
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2078_out1 = bnn_N_Mux_2_2_3_1_2077_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2078_out1 = bnn_N_Mux_2_2_3_1_2078_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2079_in1 = {s_reg_1093_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2079
         assign bnn_RightShift_64Sx8S_1S_1_2079_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2079_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2080_in3 = {bnn_RightShift_64Sx8S_1S_1_2079_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_992 or bnn_N_Mux_2_2_3_1_2080_in3)
          begin :bnn_N_Mux_2_2_3_1_2080
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2080_out1 = s_reg_992;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2080_out1 = bnn_N_Mux_2_2_3_1_2080_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_969 or s_reg_977 or s_reg_993 or bnn_N_Mux_2_2_3_1_2080_out1)
          begin :bnn_N_Mux_2_4_8_1_2081
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2081_out1 = bnn_N_Mux_2_2_3_1_2080_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2081_out1 = s_reg_993;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2081_out1 = s_reg_969;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2081_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2081_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2082
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2082_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2082_out1 = bnn_N_Mux_2_4_8_1_2081_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2083_in3 = {bnn_RightShift_64Sx8S_1S_1_1719_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2082_out1 or bnn_N_Mux_2_2_3_1_2083_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2083
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2083_out1 = bnn_N_Mux_2_2_3_1_2082_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2083_out1 = bnn_N_Mux_2_2_3_1_2083_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2084_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[20], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1968_out1 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_N_Mux_2_4_8_1_2084_in3)
          begin :bnn_N_Mux_2_4_8_1_2084
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2084_out1 = bnn_N_Mux_2_2_3_1_1968_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2084_out1 = bnn_N_Mux_2_4_8_1_2084_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2084_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2084_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2084_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2085
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2085_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2085_out1 = bnn_N_Mux_2_4_8_1_2084_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2086_in3 = {bnn_RightShift_64Sx8S_1S_1_1743_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2085_out1 or bnn_N_Mux_2_2_3_1_2086_in3)
          begin :bnn_N_Mux_2_2_3_1_2086
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2086_out1 = bnn_N_Mux_2_2_3_1_2085_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2086_out1 = bnn_N_Mux_2_2_3_1_2086_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_N_Mux_2_4_8_1_2084_in3 or bnn_N_Mux_2_2_3_1_2086_out1)
          begin :bnn_N_Mux_2_4_8_1_2087
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2087_out1 = bnn_N_Mux_2_2_3_1_2086_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2087_out1 = bnn_N_Mux_2_4_8_1_2084_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2087_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2087_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2087_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2088
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2088_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2088_out1 = bnn_N_Mux_2_4_8_1_2087_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2089_in3 = {bnn_RightShift_64Sx8S_1S_1_1663_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2088_out1 or bnn_N_Mux_2_2_3_1_2089_in3)
          begin :bnn_N_Mux_2_2_3_1_2089
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2089_out1 = bnn_N_Mux_2_2_3_1_2088_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2089_out1 = bnn_N_Mux_2_2_3_1_2089_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2090_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[28], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2080_out1 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_N_Mux_2_4_8_1_2090_in3)
          begin :bnn_N_Mux_2_4_8_1_2090
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2090_out1 = bnn_N_Mux_2_2_3_1_2080_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2090_out1 = bnn_N_Mux_2_4_8_1_2090_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2090_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2090_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2090_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2091
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2091_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2091_out1 = bnn_N_Mux_2_4_8_1_2090_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2092_in3 = {bnn_RightShift_64Sx8S_1S_1_1751_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2091_out1 or bnn_N_Mux_2_2_3_1_2092_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2092
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2092_out1 = bnn_N_Mux_2_2_3_1_2091_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2092_out1 = bnn_N_Mux_2_2_3_1_2092_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_N_Mux_2_4_8_1_2090_in3 or bnn_N_Mux_2_2_3_1_2092_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2093
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2093_out1 = bnn_N_Mux_2_2_3_1_2092_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2093_out1 = bnn_N_Mux_2_4_8_1_2090_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2093_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2093_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2093_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2094
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2094_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2094_out1 = bnn_N_Mux_2_4_8_1_2093_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2095_in3 = {bnn_RightShift_64Sx8S_1S_1_1671_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2094_out1 or bnn_N_Mux_2_2_3_1_2095_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2095
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2095_out1 = bnn_N_Mux_2_2_3_1_2094_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2095_out1 = bnn_N_Mux_2_2_3_1_2095_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2096_in1 = {s_reg_1093_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2096
         assign bnn_RightShift_64Sx8S_1S_1_2096_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2096_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2097_in3 = {bnn_RightShift_64Sx8S_1S_1_2096_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_994 or bnn_N_Mux_2_2_3_1_2097_in3)
          begin :bnn_N_Mux_2_2_3_1_2097
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2097_out1 = s_reg_994;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2097_out1 = bnn_N_Mux_2_2_3_1_2097_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_972 or s_reg_977 or s_reg_995 or bnn_N_Mux_2_2_3_1_2097_out1)
          begin :bnn_N_Mux_2_4_8_1_2098
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2098_out1 = bnn_N_Mux_2_2_3_1_2097_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2098_out1 = s_reg_995;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2098_out1 = s_reg_972;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2098_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2098_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2099
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2099_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2099_out1 = bnn_N_Mux_2_4_8_1_2098_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2100_in3 = {bnn_RightShift_64Sx8S_1S_1_1720_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2099_out1 or bnn_N_Mux_2_2_3_1_2100_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2100
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2100_out1 = bnn_N_Mux_2_2_3_1_2099_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2100_out1 = bnn_N_Mux_2_2_3_1_2100_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2101_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[21], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1979_out1 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_N_Mux_2_4_8_1_2101_in3)
          begin :bnn_N_Mux_2_4_8_1_2101
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2101_out1 = bnn_N_Mux_2_2_3_1_1979_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2101_out1 = bnn_N_Mux_2_4_8_1_2101_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2101_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2101_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2101_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2102
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2102_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2102_out1 = bnn_N_Mux_2_4_8_1_2101_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2103_in3 = {bnn_RightShift_64Sx8S_1S_1_1744_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2102_out1 or bnn_N_Mux_2_2_3_1_2103_in3)
          begin :bnn_N_Mux_2_2_3_1_2103
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2103_out1 = bnn_N_Mux_2_2_3_1_2102_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2103_out1 = bnn_N_Mux_2_2_3_1_2103_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_N_Mux_2_4_8_1_2101_in3 or bnn_N_Mux_2_2_3_1_2103_out1)
          begin :bnn_N_Mux_2_4_8_1_2104
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2104_out1 = bnn_N_Mux_2_2_3_1_2103_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2104_out1 = bnn_N_Mux_2_4_8_1_2101_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2104_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2104_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2104_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2105
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2105_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2105_out1 = bnn_N_Mux_2_4_8_1_2104_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2106_in3 = {bnn_RightShift_64Sx8S_1S_1_1664_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2105_out1 or bnn_N_Mux_2_2_3_1_2106_in3)
          begin :bnn_N_Mux_2_2_3_1_2106
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2106_out1 = bnn_N_Mux_2_2_3_1_2105_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2106_out1 = bnn_N_Mux_2_2_3_1_2106_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2107_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[29], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2097_out1 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_N_Mux_2_4_8_1_2107_in3)
          begin :bnn_N_Mux_2_4_8_1_2107
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2107_out1 = bnn_N_Mux_2_2_3_1_2097_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2107_out1 = bnn_N_Mux_2_4_8_1_2107_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2107_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2107_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2107_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2108
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2108_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2108_out1 = bnn_N_Mux_2_4_8_1_2107_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2109_in3 = {bnn_RightShift_64Sx8S_1S_1_1752_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2108_out1 or bnn_N_Mux_2_2_3_1_2109_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2109
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2109_out1 = bnn_N_Mux_2_2_3_1_2108_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2109_out1 = bnn_N_Mux_2_2_3_1_2109_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_N_Mux_2_4_8_1_2107_in3 or bnn_N_Mux_2_2_3_1_2109_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2110
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2110_out1 = bnn_N_Mux_2_2_3_1_2109_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2110_out1 = bnn_N_Mux_2_4_8_1_2107_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2110_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2110_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2110_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2111
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2111_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2111_out1 = bnn_N_Mux_2_4_8_1_2110_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2112_in3 = {bnn_RightShift_64Sx8S_1S_1_1672_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2111_out1 or bnn_N_Mux_2_2_3_1_2112_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2112
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2112_out1 = bnn_N_Mux_2_2_3_1_2111_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2112_out1 = bnn_N_Mux_2_2_3_1_2112_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2113_in1 = {s_reg_1093_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2113
         assign bnn_RightShift_64Sx8S_1S_1_2113_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2113_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2114_in3 = {bnn_RightShift_64Sx8S_1S_1_2113_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_996 or bnn_N_Mux_2_2_3_1_2114_in3)
          begin :bnn_N_Mux_2_2_3_1_2114
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2114_out1 = s_reg_996;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2114_out1 = bnn_N_Mux_2_2_3_1_2114_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_975 or s_reg_977 or s_reg_997 or bnn_N_Mux_2_2_3_1_2114_out1)
          begin :bnn_N_Mux_2_4_8_1_2115
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2115_out1 = bnn_N_Mux_2_2_3_1_2114_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2115_out1 = s_reg_997;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2115_out1 = s_reg_975;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2115_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2115_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2116
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2116_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2116_out1 = bnn_N_Mux_2_4_8_1_2115_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2117_in3 = {bnn_RightShift_64Sx8S_1S_1_1721_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2116_out1 or bnn_N_Mux_2_2_3_1_2117_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2117
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2117_out1 = bnn_N_Mux_2_2_3_1_2116_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2117_out1 = bnn_N_Mux_2_2_3_1_2117_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2118_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[22], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1990_out1 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_N_Mux_2_4_8_1_2118_in3)
          begin :bnn_N_Mux_2_4_8_1_2118
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2118_out1 = bnn_N_Mux_2_2_3_1_1990_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2118_out1 = bnn_N_Mux_2_4_8_1_2118_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2118_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2118_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2118_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2119
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2119_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2119_out1 = bnn_N_Mux_2_4_8_1_2118_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2120_in3 = {bnn_RightShift_64Sx8S_1S_1_1745_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2119_out1 or bnn_N_Mux_2_2_3_1_2120_in3)
          begin :bnn_N_Mux_2_2_3_1_2120
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2120_out1 = bnn_N_Mux_2_2_3_1_2119_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2120_out1 = bnn_N_Mux_2_2_3_1_2120_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_N_Mux_2_4_8_1_2118_in3 or bnn_N_Mux_2_2_3_1_2120_out1)
          begin :bnn_N_Mux_2_4_8_1_2121
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2121_out1 = bnn_N_Mux_2_2_3_1_2120_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2121_out1 = bnn_N_Mux_2_4_8_1_2118_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2121_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2121_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2121_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2122
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2122_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2122_out1 = bnn_N_Mux_2_4_8_1_2121_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2123_in3 = {bnn_RightShift_64Sx8S_1S_1_1665_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2122_out1 or bnn_N_Mux_2_2_3_1_2123_in3)
          begin :bnn_N_Mux_2_2_3_1_2123
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2123_out1 = bnn_N_Mux_2_2_3_1_2122_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2123_out1 = bnn_N_Mux_2_2_3_1_2123_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2124_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[30], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_2_3_1_2114_out1 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_N_Mux_2_4_8_1_2124_in3)
          begin :bnn_N_Mux_2_4_8_1_2124
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2124_out1 = bnn_N_Mux_2_2_3_1_2114_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2124_out1 = bnn_N_Mux_2_4_8_1_2124_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2124_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2124_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2124_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2125
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2125_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2125_out1 = bnn_N_Mux_2_4_8_1_2124_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2126_in3 = {bnn_RightShift_64Sx8S_1S_1_1753_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2125_out1 or bnn_N_Mux_2_2_3_1_2126_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_1_2126
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2126_out1 = bnn_N_Mux_2_2_3_1_2125_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2126_out1 = bnn_N_Mux_2_2_3_1_2126_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_N_Mux_2_4_8_1_2124_in3 or bnn_N_Mux_2_2_3_1_2126_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2127
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2127_out1 = bnn_N_Mux_2_2_3_1_2126_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2127_out1 = bnn_N_Mux_2_4_8_1_2124_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2127_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2127_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2127_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2128
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2128_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2128_out1 = bnn_N_Mux_2_4_8_1_2127_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2129_in3 = {bnn_RightShift_64Sx8S_1S_1_1673_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2128_out1 or bnn_N_Mux_2_2_3_1_2129_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_1_2129
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2129_out1 = bnn_N_Mux_2_2_3_1_2128_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2129_out1 = bnn_N_Mux_2_2_3_1_2129_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2130_in1 = {s_reg_1093_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2130
         assign bnn_RightShift_64Sx8S_1S_1_2130_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2130_in1[5:0];

         assign bnn_N_Mux_2_2_3_1_2131_in3 = {bnn_RightShift_64Sx8S_1S_1_2130_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_998 or bnn_N_Mux_2_2_3_1_2131_in3)
          begin :bnn_N_Mux_2_2_3_1_2131
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2131_out1 = s_reg_998;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2131_out1 = bnn_N_Mux_2_2_3_1_2131_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_883 or s_reg_980 or s_reg_999 or bnn_N_Mux_2_2_3_1_2131_out1)
          begin :bnn_N_Mux_2_4_8_1_2132
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2132_out1 = bnn_N_Mux_2_2_3_1_2131_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2132_out1 = s_reg_999;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2132_out1 = s_reg_980;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2132_out1 = s_reg_883;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2132_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2133
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2133_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2133_out1 = bnn_N_Mux_2_4_8_1_2132_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2134_in3 = {bnn_RightShift_64Sx8S_1S_1_1722_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2133_out1 or bnn_N_Mux_2_2_3_1_2134_in3 or s_reg_1055_stage1)
          begin :bnn_N_Mux_2_2_3_1_2134
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2134_out1 = bnn_N_Mux_2_2_3_1_2133_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2134_out1 = bnn_N_Mux_2_2_3_1_2134_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_1_2135_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[23], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2001_out1 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_N_Mux_2_4_8_1_2135_in3)
          begin :bnn_N_Mux_2_4_8_1_2135
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2135_out1 = bnn_N_Mux_2_2_3_1_2001_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2135_out1 = bnn_N_Mux_2_4_8_1_2135_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2135_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2135_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2135_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2136
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2136_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2136_out1 = bnn_N_Mux_2_4_8_1_2135_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2137_in3 = {bnn_RightShift_64Sx8S_1S_1_1746_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2136_out1 or bnn_N_Mux_2_2_3_1_2137_in3)
          begin :bnn_N_Mux_2_2_3_1_2137
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2137_out1 = bnn_N_Mux_2_2_3_1_2136_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2137_out1 = bnn_N_Mux_2_2_3_1_2137_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_N_Mux_2_4_8_1_2135_in3 or bnn_N_Mux_2_2_3_1_2137_out1)
          begin :bnn_N_Mux_2_4_8_1_2138
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2138_out1 = bnn_N_Mux_2_2_3_1_2137_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2138_out1 = bnn_N_Mux_2_4_8_1_2135_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2138_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2138_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2138_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2139
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2139_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2139_out1 = bnn_N_Mux_2_4_8_1_2138_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_2140_in3 = {bnn_RightShift_64Sx8S_1S_1_1666_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2139_out1 or bnn_N_Mux_2_2_3_1_2140_in3)
          begin :bnn_N_Mux_2_2_3_1_2140
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2140_out1 = bnn_N_Mux_2_2_3_1_2139_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2140_out1 = bnn_N_Mux_2_2_3_1_2140_in3;
            end
         end

         assign bnn_N_Mux_2_4_8_4_2141_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[31], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or s_reg_883 or bnn_N_Mux_2_2_3_1_2131_out1 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_N_Mux_2_4_8_4_2141_in3)
          begin :bnn_N_Mux_2_4_8_4_2141
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_2141_out1 = bnn_N_Mux_2_2_3_1_2131_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_2141_out1 = bnn_N_Mux_2_4_8_4_2141_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_2141_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_2141_out1 = s_reg_883;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_2141_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_4_2142
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_4_2142_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2142_out1 = bnn_N_Mux_2_4_8_4_2141_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_2143_in3 = {bnn_RightShift_64Sx8S_1S_4_1754_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_2142_out1 or bnn_N_Mux_2_2_3_4_2143_in3 or s_reg_1062_stage1)
          begin :bnn_N_Mux_2_2_3_4_2143
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_4_2143_out1 = bnn_N_Mux_2_2_3_4_2142_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2143_out1 = bnn_N_Mux_2_2_3_4_2143_in3;
            end
         end

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_N_Mux_2_4_8_4_2141_in3 or bnn_N_Mux_2_2_3_4_2143_out1 or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_2144
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_2144_out1 = bnn_N_Mux_2_2_3_4_2143_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_2144_out1 = bnn_N_Mux_2_4_8_4_2141_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_2144_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_2144_out1 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_2144_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_4_2145
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_4_2145_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2145_out1 = bnn_N_Mux_2_4_8_4_2144_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_2146_in3 = {bnn_RightShift_64Sx8S_1S_4_1674_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_2145_out1 or bnn_N_Mux_2_2_3_4_2146_in3 or s_reg_1065_stage1)
          begin :bnn_N_Mux_2_2_3_4_2146
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_4_2146_out1 = bnn_N_Mux_2_2_3_4_2145_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2146_out1 = bnn_N_Mux_2_2_3_4_2146_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2147_in1 = {s_reg_1025[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2147
         assign bnn_RightShift_64Sx8S_1S_1_2147_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2147_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_2148_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_2147_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_2148_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_2148
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_2148_out1_slice = bnn_N_Mux_3_2_6_1_2148_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_2148_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_927 or s_reg_1069_stage1 or bnn_N_Mux_3_2_6_1_2148_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2149
            if (s_reg_1069_stage1) begin
               bnn_N_Mux_2_2_3_1_2149_out1 = s_reg_927;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2149_out1 = bnn_N_Mux_3_2_6_1_2148_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_933 or s_reg_934 or s_reg_935 or bnn_N_Mux_2_2_3_1_2149_out1)
          begin :bnn_N_Mux_2_4_8_1_2150
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2150_out1 = bnn_N_Mux_2_2_3_1_2149_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2150_out1 = s_reg_934;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2150_out1 = s_reg_933;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2150_out1 = s_reg_935;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_OrReduction_10U_1U_4_1582_out1 or bnn_N_Mux_2_4_8_1_2150_out1)
          begin :bnn_N_Mux_3_2_6_1_2151
            if (bnn_OrReduction_10U_1U_4_1582_out1) begin
               bnn_N_Mux_3_2_6_1_2151_out1_slice = bnn_N_Mux_2_4_8_1_2150_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_1_2151_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1071 or bnn_N_Mux_3_2_6_1_1756_out1_slice or bnn_N_Mux_3_2_6_1_2151_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2152
            if (s_reg_1071) begin
               bnn_N_Mux_2_2_3_1_2152_out1 = bnn_N_Mux_3_2_6_1_2151_out1_slice;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2152_out1 = bnn_N_Mux_3_2_6_1_1756_out1_slice;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2153_in1 = {s_reg_886[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2153
         assign bnn_RightShift_64Sx8S_1S_1_2153_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2153_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_2154_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_2153_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_2154_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_2154
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_2154_out1_slice = bnn_N_Mux_3_2_6_1_2154_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_2154_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1077 or s_reg_946 or bnn_N_Mux_3_2_6_1_2154_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2155
            if (s_reg_1077) begin
               bnn_N_Mux_2_2_3_1_2155_out1 = s_reg_946;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2155_out1 = bnn_N_Mux_3_2_6_1_2154_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_935 or s_reg_952 or s_reg_953 or bnn_N_Mux_2_2_3_1_2155_out1)
          begin :bnn_N_Mux_2_4_8_1_2156
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2156_out1 = bnn_N_Mux_2_2_3_1_2155_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2156_out1 = s_reg_952;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2156_out1 = s_reg_935;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2156_out1 = s_reg_953;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2156_out1 or s_reg_1060_stage1)
          begin :bnn_N_Mux_2_2_3_1_2157
            if (s_reg_1060_stage1) begin
               bnn_N_Mux_2_2_3_1_2157_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2157_out1 = bnn_N_Mux_2_4_8_1_2156_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2157_out1 or s_reg_1049_stage1 or bnn_N_Mux_3_2_6_1_1758_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2158
            if (s_reg_1049_stage1) begin
               bnn_N_Mux_2_2_3_1_2158_out1 = bnn_N_Mux_2_2_3_1_2157_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2158_out1 = bnn_N_Mux_3_2_6_1_1758_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_1928_in3 or bnn_N_Mux_2_2_3_1_2149_out1 or bnn_N_Mux_2_2_3_1_2152_out1 or bnn_N_Mux_2_2_3_1_2158_out1)
          begin :bnn_N_Mux_2_4_8_1_2159
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2159_out1 = bnn_N_Mux_2_2_3_1_2149_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2159_out1 = bnn_N_Mux_2_4_8_1_1928_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2159_out1 = bnn_N_Mux_2_2_3_1_2152_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2159_out1 = bnn_N_Mux_2_2_3_1_2158_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2159_out1 or s_reg_1050_stage1)
          begin :bnn_N_Mux_2_2_3_1_2160
            if (s_reg_1050_stage1) begin
               bnn_N_Mux_2_2_3_1_2160_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2160_out1 = bnn_N_Mux_2_4_8_1_2159_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2160_out1 or s_reg_1037_stage1 or bnn_N_Mux_3_2_6_1_1766_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2161
            if (s_reg_1037_stage1) begin
               bnn_N_Mux_2_2_3_1_2161_out1 = bnn_N_Mux_2_2_3_1_2160_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2161_out1 = bnn_N_Mux_3_2_6_1_1766_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_1928_in3 or bnn_N_Mux_2_2_3_1_2152_out1 or bnn_N_Mux_2_2_3_1_2158_out1 or bnn_N_Mux_2_2_3_1_2161_out1)
          begin :bnn_N_Mux_2_4_8_1_2162
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2162_out1 = bnn_N_Mux_2_2_3_1_2161_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2162_out1 = bnn_N_Mux_2_4_8_1_1928_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2162_out1 = bnn_N_Mux_2_2_3_1_2152_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2162_out1 = bnn_N_Mux_2_2_3_1_2158_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2162_out1 or s_reg_1053_stage1)
          begin :bnn_N_Mux_2_2_3_1_2163
            if (s_reg_1053_stage1) begin
               bnn_N_Mux_2_2_3_1_2163_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2163_out1 = bnn_N_Mux_2_4_8_1_2162_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2163_out1 or s_reg_1038_stage1 or bnn_N_Mux_3_2_6_1_1676_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2164
            if (s_reg_1038_stage1) begin
               bnn_N_Mux_2_2_3_1_2164_out1 = bnn_N_Mux_2_2_3_1_2163_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2164_out1 = bnn_N_Mux_3_2_6_1_1676_out1_slice;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2165
         assign bnn_RightShift_64Sx8S_1S_1_2165_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1089[5:0];

         assign bnn_N_Mux_3_2_6_1_2166_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_2165_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_2166_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_2166
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_2166_out1_slice = bnn_N_Mux_3_2_6_1_2166_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_2166_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_943 or bnn_N_Mux_3_2_6_1_2166_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2167
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_2167_out1 = s_reg_943;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2167_out1 = bnn_N_Mux_3_2_6_1_2166_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_905 or s_reg_948 or s_reg_950 or bnn_N_Mux_2_2_3_1_2167_out1)
          begin :bnn_N_Mux_2_4_8_1_2168
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2168_out1 = bnn_N_Mux_2_2_3_1_2167_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2168_out1 = s_reg_948;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2168_out1 = s_reg_905;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2168_out1 = s_reg_950;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2168_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_2169
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_2169_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2169_out1 = bnn_N_Mux_2_4_8_1_2168_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_2169_out1 or bnn_N_Mux_3_2_6_1_1760_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2170
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_2170_out1 = bnn_N_Mux_2_2_3_1_2169_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2170_out1 = bnn_N_Mux_3_2_6_1_1760_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_1907_in3 or bnn_N_Mux_2_2_3_1_1915_out1 or bnn_N_Mux_2_2_3_1_1918_out1 or bnn_N_Mux_2_2_3_1_2170_out1)
          begin :bnn_N_Mux_2_4_8_1_2171
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2171_out1 = bnn_N_Mux_2_2_3_1_1915_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2171_out1 = bnn_N_Mux_2_4_8_1_1907_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2171_out1 = bnn_N_Mux_2_2_3_1_1918_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2171_out1 = bnn_N_Mux_2_2_3_1_2170_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2171_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_2172
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_2172_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2172_out1 = bnn_N_Mux_2_4_8_1_2171_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2172_out1 or s_reg_1051_stage1 or bnn_N_Mux_3_2_6_1_1768_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2173
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_2173_out1 = bnn_N_Mux_2_2_3_1_2172_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2173_out1 = bnn_N_Mux_3_2_6_1_1768_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_1907_in3 or bnn_N_Mux_2_2_3_1_1918_out1 or bnn_N_Mux_2_2_3_1_2170_out1 or bnn_N_Mux_2_2_3_1_2173_out1)
          begin :bnn_N_Mux_2_4_8_1_2174
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2174_out1 = bnn_N_Mux_2_2_3_1_2173_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2174_out1 = bnn_N_Mux_2_4_8_1_1907_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2174_out1 = bnn_N_Mux_2_2_3_1_1918_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2174_out1 = bnn_N_Mux_2_2_3_1_2170_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2174_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_2175
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_2175_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2175_out1 = bnn_N_Mux_2_4_8_1_2174_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_2175_out1 or bnn_N_Mux_3_2_6_1_1678_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2176
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_2176_out1 = bnn_N_Mux_2_2_3_1_2175_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2176_out1 = bnn_N_Mux_3_2_6_1_1678_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_7_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2176_out1 or bnn_N_Mux_3_2_6_4_1920_out1_slice or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :bnn_N_Mux_2_4_7_4_2177
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_7_4_2177_out1 = bnn_N_Mux_3_2_6_4_1920_out1_slice;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_7_4_2177_out1 = 2'd0;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_7_4_2177_out1 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
               end
               
               default: begin
                  bnn_N_Mux_2_4_7_4_2177_out1 = bnn_N_Mux_2_2_3_1_2176_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_And_1Sx1U_1U_4_1580_out1 or bnn_N_Mux_2_4_7_4_2177_out1)
          begin :bnn_N_Mux_3_2_6_4_2178
            if (bnn_And_1Sx1U_1U_4_1580_out1) begin
               bnn_N_Mux_3_2_6_4_2178_out1_slice = bnn_N_Mux_2_4_7_4_2177_out1;
            end
            else begin
               bnn_N_Mux_3_2_6_4_2178_out1_slice = 2'd0;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_2179_in1 = {s_reg_1097[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2179
         assign bnn_RightShift_64Sx8S_1S_1_2179_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_2179_in1[5:0];

         assign bnn_N_Mux_3_2_6_1_2180_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_2179_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_2180_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_2180
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_2180_out1_slice = bnn_N_Mux_3_2_6_1_2180_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_2180_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1087 or s_reg_979 or bnn_N_Mux_3_2_6_1_2180_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2181
            if (s_reg_1087) begin
               bnn_N_Mux_2_2_3_1_2181_out1 = s_reg_979;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2181_out1 = bnn_N_Mux_3_2_6_1_2180_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_953 or s_reg_983 or s_reg_984 or bnn_N_Mux_2_2_3_1_2181_out1)
          begin :bnn_N_Mux_2_4_8_1_2182
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2182_out1 = bnn_N_Mux_2_2_3_1_2181_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2182_out1 = s_reg_983;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2182_out1 = s_reg_953;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2182_out1 = s_reg_984;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2182_out1 or s_reg_1085_stage1)
          begin :bnn_N_Mux_2_2_3_1_2183
            if (s_reg_1085_stage1) begin
               bnn_N_Mux_2_2_3_1_2183_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2183_out1 = bnn_N_Mux_2_4_8_1_2182_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1084 or bnn_N_Mux_2_2_3_1_2183_out1 or bnn_N_Mux_3_2_6_1_1762_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2184
            if (s_reg_1084) begin
               bnn_N_Mux_2_2_3_1_2184_out1 = bnn_N_Mux_2_2_3_1_2183_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2184_out1 = bnn_N_Mux_3_2_6_1_1762_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2155_out1 or bnn_N_Mux_2_2_3_1_2158_out1 or bnn_N_Mux_2_2_3_1_2184_out1 or bnn_N_Mux_3_2_6_1_1687_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2185
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2185_out1 = bnn_N_Mux_2_2_3_1_2155_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2185_out1 = bnn_N_Mux_3_2_6_1_1687_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2185_out1 = bnn_N_Mux_2_2_3_1_2158_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2185_out1 = bnn_N_Mux_2_2_3_1_2184_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2185_out1 or s_reg_1052_stage1)
          begin :bnn_N_Mux_2_2_3_1_2186
            if (s_reg_1052_stage1) begin
               bnn_N_Mux_2_2_3_1_2186_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2186_out1 = bnn_N_Mux_2_4_8_1_2185_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2186_out1 or s_reg_1051_stage1 or bnn_N_Mux_3_2_6_1_1770_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2187
            if (s_reg_1051_stage1) begin
               bnn_N_Mux_2_2_3_1_2187_out1 = bnn_N_Mux_2_2_3_1_2186_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2187_out1 = bnn_N_Mux_3_2_6_1_1770_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2158_out1 or bnn_N_Mux_2_2_3_1_2184_out1 or bnn_N_Mux_2_2_3_1_2187_out1 or bnn_N_Mux_3_2_6_1_1687_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2188
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2188_out1 = bnn_N_Mux_2_2_3_1_2187_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2188_out1 = bnn_N_Mux_3_2_6_1_1687_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2188_out1 = bnn_N_Mux_2_2_3_1_2158_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2188_out1 = bnn_N_Mux_2_2_3_1_2184_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2188_out1 or s_reg_1054_stage1)
          begin :bnn_N_Mux_2_2_3_1_2189
            if (s_reg_1054_stage1) begin
               bnn_N_Mux_2_2_3_1_2189_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2189_out1 = bnn_N_Mux_2_4_8_1_2188_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1579_out1 or bnn_N_Mux_2_2_3_1_2189_out1 or bnn_N_Mux_3_2_6_1_1680_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2190
            if (bnn_Or_1Sx1U_1S_4_1579_out1) begin
               bnn_N_Mux_2_2_3_1_2190_out1 = bnn_N_Mux_2_2_3_1_2189_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2190_out1 = bnn_N_Mux_3_2_6_1_1680_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_2022_in3 or bnn_N_Mux_2_2_3_1_2181_out1 or bnn_N_Mux_2_2_3_1_2184_out1 or bnn_N_Mux_3_2_6_1_1783_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2191
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2191_out1 = bnn_N_Mux_2_2_3_1_2181_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2191_out1 = bnn_N_Mux_2_4_8_1_2022_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2191_out1 = bnn_N_Mux_2_2_3_1_2184_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2191_out1 = bnn_N_Mux_3_2_6_1_1783_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2191_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2192
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2192_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2192_out1 = bnn_N_Mux_2_4_8_1_2191_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2192_out1 or bnn_N_Mux_3_2_6_1_1774_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2193
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2193_out1 = bnn_N_Mux_2_2_3_1_2192_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2193_out1 = bnn_N_Mux_3_2_6_1_1774_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_2022_in3 or bnn_N_Mux_2_2_3_1_2184_out1 or bnn_N_Mux_2_2_3_1_2193_out1 or bnn_N_Mux_3_2_6_1_1783_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2194
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2194_out1 = bnn_N_Mux_2_2_3_1_2193_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2194_out1 = bnn_N_Mux_2_4_8_1_2022_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2194_out1 = bnn_N_Mux_2_2_3_1_2184_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2194_out1 = bnn_N_Mux_3_2_6_1_1783_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2194_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2195
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2195_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2195_out1 = bnn_N_Mux_2_4_8_1_2194_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2195_out1 or bnn_N_Mux_3_2_6_1_1684_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2196
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2196_out1 = bnn_N_Mux_2_2_3_1_2195_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2196_out1 = bnn_N_Mux_3_2_6_1_1684_out1_slice;
            end
         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_2197
         assign bnn_RightShift_64Sx8S_1S_1_2197_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> s_reg_1096[5:0];

         assign bnn_N_Mux_3_2_6_1_2198_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_2197_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_2198_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_2198
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_2198_out1_slice = bnn_N_Mux_3_2_6_1_2198_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_2198_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1094 or s_reg_976 or bnn_N_Mux_3_2_6_1_2198_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2199
            if (s_reg_1094) begin
               bnn_N_Mux_2_2_3_1_2199_out1 = s_reg_976;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2199_out1 = bnn_N_Mux_3_2_6_1_2198_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_950 or s_reg_977 or s_reg_981 or bnn_N_Mux_2_2_3_1_2199_out1)
          begin :bnn_N_Mux_2_4_8_1_2200
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2200_out1 = bnn_N_Mux_2_2_3_1_2199_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2200_out1 = s_reg_981;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2200_out1 = s_reg_950;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2200_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2200_out1 or s_reg_1079_stage1)
          begin :bnn_N_Mux_2_2_3_1_2201
            if (s_reg_1079_stage1) begin
               bnn_N_Mux_2_2_3_1_2201_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2201_out1 = bnn_N_Mux_2_4_8_1_2200_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2201_out1 or s_reg_1055_stage1 or bnn_N_Mux_3_2_6_1_1764_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2202
            if (s_reg_1055_stage1) begin
               bnn_N_Mux_2_2_3_1_2202_out1 = bnn_N_Mux_2_2_3_1_2201_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2202_out1 = bnn_N_Mux_3_2_6_1_1764_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2167_out1 or bnn_N_Mux_2_2_3_1_2170_out1 or bnn_N_Mux_2_2_3_1_2202_out1 or bnn_N_Mux_3_2_6_1_1688_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2203
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2203_out1 = bnn_N_Mux_2_2_3_1_2167_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2203_out1 = bnn_N_Mux_3_2_6_1_1688_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2203_out1 = bnn_N_Mux_2_2_3_1_2170_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2203_out1 = bnn_N_Mux_2_2_3_1_2202_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2203_out1 or s_reg_1073_stage1)
          begin :bnn_N_Mux_2_2_3_1_2204
            if (s_reg_1073_stage1) begin
               bnn_N_Mux_2_2_3_1_2204_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2204_out1 = bnn_N_Mux_2_4_8_1_2203_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_1072 or bnn_N_Mux_2_2_3_1_2204_out1 or bnn_N_Mux_3_2_6_1_1772_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2205
            if (s_reg_1072) begin
               bnn_N_Mux_2_2_3_1_2205_out1 = bnn_N_Mux_2_2_3_1_2204_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2205_out1 = bnn_N_Mux_3_2_6_1_1772_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2170_out1 or bnn_N_Mux_2_2_3_1_2202_out1 or bnn_N_Mux_2_2_3_1_2205_out1 or bnn_N_Mux_3_2_6_1_1688_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2206
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2206_out1 = bnn_N_Mux_2_2_3_1_2205_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2206_out1 = bnn_N_Mux_3_2_6_1_1688_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2206_out1 = bnn_N_Mux_2_2_3_1_2170_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2206_out1 = bnn_N_Mux_2_2_3_1_2202_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2206_out1 or s_reg_1074_stage1)
          begin :bnn_N_Mux_2_2_3_1_2207
            if (s_reg_1074_stage1) begin
               bnn_N_Mux_2_2_3_1_2207_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2207_out1 = bnn_N_Mux_2_4_8_1_2206_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1586_out1 or bnn_N_Mux_2_2_3_1_2207_out1 or bnn_N_Mux_3_2_6_1_1682_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2208
            if (bnn_Or_1Sx1U_1S_4_1586_out1) begin
               bnn_N_Mux_2_2_3_1_2208_out1 = bnn_N_Mux_2_2_3_1_2207_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2208_out1 = bnn_N_Mux_3_2_6_1_1682_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or s_reg_977 or bnn_N_Mux_2_4_8_1_2135_in3 or bnn_N_Mux_2_2_3_1_2199_out1 or bnn_N_Mux_2_2_3_1_2202_out1)
          begin :bnn_N_Mux_2_4_8_1_2209
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2209_out1 = bnn_N_Mux_2_2_3_1_2199_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2209_out1 = bnn_N_Mux_2_4_8_1_2135_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2209_out1 = bnn_N_Mux_2_2_3_1_2202_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2209_out1 = s_reg_977;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2209_out1 or s_reg_1080_stage1)
          begin :bnn_N_Mux_2_2_3_1_2210
            if (s_reg_1080_stage1) begin
               bnn_N_Mux_2_2_3_1_2210_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2210_out1 = bnn_N_Mux_2_4_8_1_2209_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2210_out1 or s_reg_1062_stage1 or bnn_N_Mux_3_2_6_1_1776_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2211
            if (s_reg_1062_stage1) begin
               bnn_N_Mux_2_2_3_1_2211_out1 = bnn_N_Mux_2_2_3_1_2210_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2211_out1 = bnn_N_Mux_3_2_6_1_1776_out1_slice;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_4_8_1_2135_in3 or bnn_N_Mux_2_2_3_1_2202_out1 or bnn_N_Mux_2_2_3_1_2211_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_2212
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_2212_out1 = bnn_N_Mux_2_2_3_1_2211_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_2212_out1 = bnn_N_Mux_2_4_8_1_2135_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_2212_out1 = bnn_N_Mux_2_2_3_1_2202_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_2212_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_2212_out1 or s_reg_1081_stage1)
          begin :bnn_N_Mux_2_2_3_1_2213
            if (s_reg_1081_stage1) begin
               bnn_N_Mux_2_2_3_1_2213_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2213_out1 = bnn_N_Mux_2_4_8_1_2212_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_2213_out1 or s_reg_1065_stage1 or bnn_N_Mux_3_2_6_1_1686_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_2214
            if (s_reg_1065_stage1) begin
               bnn_N_Mux_2_2_3_1_2214_out1 = bnn_N_Mux_2_2_3_1_2213_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2214_out1 = bnn_N_Mux_3_2_6_1_1686_out1_slice;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2215
         assign bnn_Minus_2S_2S_1_2215_out1 = -bnn_N_Mux_2_2_3_1_1790_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2216
         assign bnn_Minus_2S_2S_1_2216_out1 = -bnn_N_Mux_2_2_3_1_1781_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1790_out1 or bnn_Minus_2S_2S_1_2215_out1)
          begin :bnn_N_Mux_2_2_3_1_2218
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2218_out1 = bnn_Minus_2S_2S_1_2215_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2218_out1 = bnn_N_Mux_2_2_3_1_1790_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1781_out1 or bnn_Minus_2S_2S_1_2216_out1)
          begin :bnn_N_Mux_2_2_3_1_2219
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2219_out1 = bnn_Minus_2S_2S_1_2216_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2219_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2220
         assign bnn_Minus_2S_2S_1_2220_out1 = -bnn_N_Mux_2_2_3_1_1795_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1781_out1 or bnn_Minus_2S_2S_1_2216_out1)
          begin :bnn_N_Mux_2_2_3_1_2223
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2223_out1 = bnn_Minus_2S_2S_1_2216_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2223_out1 = bnn_N_Mux_2_2_3_1_1781_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2225
         assign bnn_Minus_2S_2S_1_2225_out1 = -bnn_N_Mux_2_4_8_1_1826_in3;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2226
         assign bnn_Add_2Sx2S_3S_1_2226_out1 = {bnn_N_Mux_2_2_3_1_2219_out1[1], bnn_N_Mux_2_2_3_1_2219_out1} + {bnn_N_Mux_2_2_3_1_2218_out1[1], bnn_N_Mux_2_2_3_1_2218_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1795_out1 or bnn_Minus_2S_2S_1_2220_out1)
          begin :bnn_N_Mux_2_2_3_1_2227
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_2227_out1 = bnn_Minus_2S_2S_1_2220_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2227_out1 = bnn_N_Mux_2_2_3_1_1795_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1795_out1 or bnn_Minus_2S_2S_1_2220_out1)
          begin :bnn_N_Mux_2_2_3_1_2228
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2228_out1 = bnn_Minus_2S_2S_1_2220_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2228_out1 = bnn_N_Mux_2_2_3_1_1795_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1790_out1 or bnn_Minus_2S_2S_1_2215_out1)
          begin :bnn_N_Mux_2_2_3_1_2229
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2229_out1 = bnn_Minus_2S_2S_1_2215_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2229_out1 = bnn_N_Mux_2_2_3_1_1790_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2230
         assign bnn_Minus_2S_2S_1_2230_out1 = -bnn_N_Mux_2_2_3_1_1800_out1;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2234
         assign bnn_Add_2Sx2S_3S_1_2234_out1 = {bnn_N_Mux_2_2_3_4_1634_out1[1], bnn_N_Mux_2_2_3_4_1634_out1} + {bnn_N_Mux_2_2_3_1_2223_out1[1], bnn_N_Mux_2_2_3_1_2223_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1790_out1 or bnn_Minus_2S_2S_1_2215_out1)
          begin :bnn_N_Mux_2_2_3_1_2235
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_2235_out1 = bnn_Minus_2S_2S_1_2215_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2235_out1 = bnn_N_Mux_2_2_3_1_1790_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2236
         assign bnn_Minus_2S_2S_1_2236_out1 = -bnn_N_Mux_2_4_8_1_1841_in3;

         assign bnn_N_Mux_2_2_3_1_2237_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[0], 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_2225_out1 or bnn_N_Mux_2_2_3_1_2237_in3)
          begin :bnn_N_Mux_2_2_3_1_2237
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_2237_out1 = bnn_Minus_2S_2S_1_2225_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2237_out1 = bnn_N_Mux_2_2_3_1_2237_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2238
         assign bnn_Add_3Sx3S_4S_1_2238_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_2227_out1[1]}}, bnn_N_Mux_2_2_3_1_2227_out1} + {bnn_Add_2Sx2S_3S_1_2226_out1[2], bnn_Add_2Sx2S_3S_1_2226_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2240
         assign bnn_Add_2Sx2S_3S_1_2240_out1 = {bnn_N_Mux_2_2_3_1_2229_out1[1], bnn_N_Mux_2_2_3_1_2229_out1} + {bnn_N_Mux_2_2_3_1_2228_out1[1], bnn_N_Mux_2_2_3_1_2228_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1800_out1 or bnn_Minus_2S_2S_1_2230_out1)
          begin :bnn_N_Mux_2_2_3_1_2241
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_2241_out1 = bnn_Minus_2S_2S_1_2230_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2241_out1 = bnn_N_Mux_2_2_3_1_1800_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1800_out1 or bnn_Minus_2S_2S_1_2230_out1)
          begin :bnn_N_Mux_2_2_3_1_2242
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2242_out1 = bnn_Minus_2S_2S_1_2230_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2242_out1 = bnn_N_Mux_2_2_3_1_1800_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1795_out1 or bnn_Minus_2S_2S_1_2220_out1)
          begin :bnn_N_Mux_2_2_3_1_2243
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2243_out1 = bnn_Minus_2S_2S_1_2220_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2243_out1 = bnn_N_Mux_2_2_3_1_1795_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_953 or bnn_N_Mux_2_2_3_1_1805_out1 or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_1_2244_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_1_2244_in1 = s_reg_953;
            end
            else begin
               bnn_Minus_2S_2S_1_2244_in1 = bnn_N_Mux_2_2_3_1_1805_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2244
         assign bnn_Minus_2S_2S_1_2244_out1 = -bnn_Minus_2S_2S_1_2244_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_1_2225_out1 or bnn_N_Mux_2_2_3_1_2237_in3)
          begin :bnn_N_Mux_2_2_3_4_2248
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2248_out1 = bnn_Minus_2S_2S_1_2225_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2248_out1 = bnn_N_Mux_2_2_3_1_2237_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2249
         assign bnn_Add_3Sx3S_4S_1_2249_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_2235_out1[1]}}, bnn_N_Mux_2_2_3_1_2235_out1} + {bnn_Add_2Sx2S_3S_1_2234_out1[2], bnn_Add_2Sx2S_3S_1_2234_out1};

         // resource: mux_2bx2i
         always @(s_reg_973 or bnn_N_Mux_64_2_2_1_1636_out1[2] or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_1_2250_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_1_2250_in1 = s_reg_973;
            end
            else begin
               bnn_Minus_2S_2S_1_2250_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[2], 1'b1};
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2250
         assign bnn_Minus_2S_2S_1_2250_out1 = -bnn_Minus_2S_2S_1_2250_in1;

         assign bnn_N_Mux_2_2_3_1_2251_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[1], 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_2236_out1 or bnn_N_Mux_2_2_3_1_2251_in3)
          begin :bnn_N_Mux_2_2_3_1_2251
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_2251_out1 = bnn_Minus_2S_2S_1_2236_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2251_out1 = bnn_N_Mux_2_2_3_1_2251_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2252
         assign bnn_Add_4Sx2S_4S_1_2252_out1 = bnn_Add_3Sx3S_4S_1_2238_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_2237_out1[1]}}, bnn_N_Mux_2_2_3_1_2237_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_2236_out1 or bnn_N_Mux_2_2_3_1_2251_in3)
          begin :bnn_N_Mux_2_2_3_1_2254
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_2254_out1 = bnn_Minus_2S_2S_1_2236_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2254_out1 = bnn_N_Mux_2_2_3_1_2251_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2255
         assign bnn_Add_3Sx3S_4S_1_2255_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_2241_out1[1]}}, bnn_N_Mux_2_2_3_1_2241_out1} + {bnn_Add_2Sx2S_3S_1_2240_out1[2], bnn_Add_2Sx2S_3S_1_2240_out1};

         // resource: mux_2bx2i
         always @(s_reg_1119[1:0] or bnn_N_Mux_2_2_3_1_2243_out1 or gs_ctrl105)
          begin :drive_bnn_Add_2Sx2S_3S_1_2257_in2
            if (gs_ctrl105) begin
               bnn_Add_2Sx2S_3S_1_2257_in2 = s_reg_1119[1:0];
            end
            else begin
               bnn_Add_2Sx2S_3S_1_2257_in2 = bnn_N_Mux_2_2_3_1_2243_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1118[1:0] or bnn_N_Mux_2_2_3_1_2242_out1 or gs_ctrl105)
          begin :drive_bnn_Add_2Sx2S_3S_1_2257_in1
            if (gs_ctrl105) begin
               bnn_Add_2Sx2S_3S_1_2257_in1 = s_reg_1118[1:0];
            end
            else begin
               bnn_Add_2Sx2S_3S_1_2257_in1 = bnn_N_Mux_2_2_3_1_2242_out1;
            end
         end

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2257
         assign bnn_Add_2Sx2S_3S_1_2257_out1 = {bnn_Add_2Sx2S_3S_1_2257_in2[1], bnn_Add_2Sx2S_3S_1_2257_in2} + {bnn_Add_2Sx2S_3S_1_2257_in1[1], bnn_Add_2Sx2S_3S_1_2257_in1};

         // resource: mux_2bx2i
         always @(s_reg_953 or bnn_N_Mux_2_2_3_1_1805_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_2258_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_2258_in3 = s_reg_953;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2258_in3 = bnn_N_Mux_2_2_3_1_1805_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_2244_out1 or bnn_N_Mux_2_2_3_1_2258_in3)
          begin :bnn_N_Mux_2_2_3_1_2258
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_2258_out1 = bnn_Minus_2S_2S_1_2244_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2258_out1 = bnn_N_Mux_2_2_3_1_2258_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1805_out1 or bnn_Minus_2S_2S_1_2244_out1)
          begin :bnn_N_Mux_2_2_3_1_2259
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2259_out1 = bnn_Minus_2S_2S_1_2244_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2259_out1 = bnn_N_Mux_2_2_3_1_1805_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1800_out1 or bnn_Minus_2S_2S_1_2230_out1)
          begin :bnn_N_Mux_2_2_3_1_2260
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2260_out1 = bnn_Minus_2S_2S_1_2230_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2260_out1 = bnn_N_Mux_2_2_3_1_1800_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2261
         assign bnn_Minus_2S_2S_1_2261_out1 = -bnn_N_Mux_2_2_3_1_1810_out1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2264
         assign bnn_Minus_2S_2S_4_2264_out1 = -bnn_N_Mux_3_2_6_4_1920_out1_slice;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_1_2236_out1 or bnn_N_Mux_2_2_3_1_2251_in3)
          begin :bnn_N_Mux_2_2_3_4_2265
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2265_out1 = bnn_Minus_2S_2S_1_2236_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2265_out1 = bnn_N_Mux_2_2_3_1_2251_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2266
         assign bnn_Add_4Sx2S_4S_1_2266_out1 = bnn_Add_3Sx3S_4S_1_2249_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2248_out1[1]}}, bnn_N_Mux_2_2_3_4_2248_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2267
         assign bnn_Minus_2S_2S_4_2267_out1 = -bnn_N_Mux_2_2_3_1_1828_out1;

         // resource: mux_2bx2i
         always @(s_reg_973 or bnn_N_Mux_64_2_2_1_1636_out1[2] or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_4_2268_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_4_2268_in3 = s_reg_973;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2268_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[2], 1'b1};
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_1_2250_out1 or bnn_N_Mux_2_2_3_4_2268_in3)
          begin :bnn_N_Mux_2_2_3_4_2268
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2268_out1 = bnn_Minus_2S_2S_1_2250_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2268_out1 = bnn_N_Mux_2_2_3_4_2268_in3;
            end
         end

         // resource: mux_4bx2i
         always @(s_reg_1028 or bnn_Add_4Sx2S_4S_1_2252_out1 or gs_ctrl105)
          begin :drive_bnn_Add_4Sx2S_4S_1_2269_in2
            if (gs_ctrl105) begin
               bnn_Add_4Sx2S_4S_1_2269_in2 = s_reg_1028;
            end
            else begin
               bnn_Add_4Sx2S_4S_1_2269_in2 = bnn_Add_4Sx2S_4S_1_2252_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1123[1:0] or bnn_N_Mux_2_2_3_1_2251_out1 or gs_ctrl105)
          begin :drive_bnn_Add_4Sx2S_4S_1_2269_in1
            if (gs_ctrl105) begin
               bnn_Add_4Sx2S_4S_1_2269_in1 = s_reg_1123[1:0];
            end
            else begin
               bnn_Add_4Sx2S_4S_1_2269_in1 = bnn_N_Mux_2_2_3_1_2251_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2269
         assign bnn_Add_4Sx2S_4S_1_2269_out1 = bnn_Add_4Sx2S_4S_1_2269_in2 + {{ 2 {bnn_Add_4Sx2S_4S_1_2269_in1[1]}}, bnn_Add_4Sx2S_4S_1_2269_in1};

         // resource: mux_2bx2i
         always @(s_reg_978 or bnn_N_Mux_64_2_2_1_1636_out1[3] or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_1_2270_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_1_2270_in1 = s_reg_978;
            end
            else begin
               bnn_Minus_2S_2S_1_2270_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[3], 1'b1};
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2270
         assign bnn_Minus_2S_2S_1_2270_out1 = -bnn_Minus_2S_2S_1_2270_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_2250_out1 or bnn_N_Mux_2_2_3_4_2268_in3)
          begin :bnn_N_Mux_2_2_3_1_2271
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_2271_out1 = bnn_Minus_2S_2S_1_2250_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2271_out1 = bnn_N_Mux_2_2_3_4_2268_in3;
            end
         end

         // resource: mux_4bx2i
         always @(s_reg_1027[3:0] or bnn_Add_3Sx3S_4S_1_2255_out1 or gs_ctrl105)
          begin :drive_bnn_Add_4Sx2S_4S_1_2272_in2
            if (gs_ctrl105) begin
               bnn_Add_4Sx2S_4S_1_2272_in2 = s_reg_1027[3:0];
            end
            else begin
               bnn_Add_4Sx2S_4S_1_2272_in2 = bnn_Add_3Sx3S_4S_1_2255_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1124[1:0] or bnn_N_Mux_2_2_3_1_2254_out1 or gs_ctrl105)
          begin :drive_bnn_Add_4Sx2S_4S_1_2272_in1
            if (gs_ctrl105) begin
               bnn_Add_4Sx2S_4S_1_2272_in1 = s_reg_1124[1:0];
            end
            else begin
               bnn_Add_4Sx2S_4S_1_2272_in1 = bnn_N_Mux_2_2_3_1_2254_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2272
         assign bnn_Add_4Sx2S_4S_1_2272_out1 = bnn_Add_4Sx2S_4S_1_2272_in2 + {{ 2 {bnn_Add_4Sx2S_4S_1_2272_in1[1]}}, bnn_Add_4Sx2S_4S_1_2272_in1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_924 or bnn_Minus_2S_2S_1_2250_out1 or bnn_N_Mux_2_2_3_4_2268_in3)
          begin :bnn_N_Mux_2_2_3_1_2274
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_1_2274_out1 = bnn_Minus_2S_2S_1_2250_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2274_out1 = bnn_N_Mux_2_2_3_4_2268_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2275
         assign bnn_Add_3Sx3S_4S_1_2275_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_2258_out1[1]}}, bnn_N_Mux_2_2_3_1_2258_out1} + {bnn_Add_2Sx2S_3S_1_2257_out1[2], bnn_Add_2Sx2S_3S_1_2257_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2277
         assign bnn_Add_2Sx2S_3S_1_2277_out1 = {bnn_N_Mux_2_2_3_1_2260_out1[1], bnn_N_Mux_2_2_3_1_2260_out1} + {bnn_N_Mux_2_2_3_1_2259_out1[1], bnn_N_Mux_2_2_3_1_2259_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1810_out1 or bnn_Minus_2S_2S_1_2261_out1)
          begin :bnn_N_Mux_2_2_3_4_2278
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2278_out1 = bnn_Minus_2S_2S_1_2261_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2278_out1 = bnn_N_Mux_2_2_3_1_1810_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1810_out1 or bnn_Minus_2S_2S_1_2261_out1)
          begin :bnn_N_Mux_2_2_3_1_2279
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2279_out1 = bnn_Minus_2S_2S_1_2261_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2279_out1 = bnn_N_Mux_2_2_3_1_1810_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1805_out1 or bnn_Minus_2S_2S_1_2244_out1)
          begin :bnn_N_Mux_2_2_3_1_2280
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2280_out1 = bnn_Minus_2S_2S_1_2244_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2280_out1 = bnn_N_Mux_2_2_3_1_1805_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2281
         assign bnn_Minus_2S_2S_1_2281_out1 = -bnn_N_Mux_2_2_3_1_1815_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_Minus_2S_2S_4_2264_out1 or bnn_N_Mux_3_2_6_4_1920_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2285
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2285_out1 = bnn_Minus_2S_2S_4_2264_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2285_out1 = bnn_N_Mux_3_2_6_4_1920_out1_slice;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2286
         assign bnn_Add_4Sx2S_4S_1_2286_out1 = bnn_Add_4Sx2S_4S_1_2266_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2265_out1[1]}}, bnn_N_Mux_2_2_3_4_2265_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2287
         assign bnn_Minus_2S_2S_4_2287_out1 = -bnn_N_Mux_2_2_3_1_1843_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1828_out1 or bnn_Minus_2S_2S_4_2267_out1)
          begin :bnn_N_Mux_2_2_3_4_2288
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2288_out1 = bnn_Minus_2S_2S_4_2267_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2288_out1 = bnn_N_Mux_2_2_3_1_1828_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2289
         assign bnn_Add_4Sx2S_5S_1_2289_out1 = {bnn_Add_4Sx2S_4S_1_2269_out1[3], bnn_Add_4Sx2S_4S_1_2269_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2268_out1[1]}}, bnn_N_Mux_2_2_3_4_2268_out1};

         // resource: mux_2bx2i
         always @(s_reg_978 or bnn_N_Mux_64_2_2_1_1636_out1[3] or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_2291_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_2291_in3 = s_reg_978;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2291_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[3], 1'b1};
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_2270_out1 or bnn_N_Mux_2_2_3_1_2291_in3)
          begin :bnn_N_Mux_2_2_3_1_2291
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_2291_out1 = bnn_Minus_2S_2S_1_2270_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2291_out1 = bnn_N_Mux_2_2_3_1_2291_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2292
         assign bnn_Add_4Sx2S_4S_1_2292_out1 = bnn_Add_4Sx2S_4S_1_2272_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_2271_out1[1]}}, bnn_N_Mux_2_2_3_1_2271_out1};

         // resource: mux_2bx2i
         always @(s_reg_983 or bnn_N_Mux_64_2_2_1_1636_out1[4] or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_1_2293_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_1_2293_in1 = s_reg_983;
            end
            else begin
               bnn_Minus_2S_2S_1_2293_in1 = {bnn_N_Mux_64_2_2_1_1636_out1[4], 1'b1};
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2293
         assign bnn_Minus_2S_2S_1_2293_out1 = -bnn_Minus_2S_2S_1_2293_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_932 or bnn_Minus_2S_2S_1_2270_out1 or bnn_N_Mux_2_2_3_1_2291_in3)
          begin :bnn_N_Mux_2_2_3_1_2294
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_1_2294_out1 = bnn_Minus_2S_2S_1_2270_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2294_out1 = bnn_N_Mux_2_2_3_1_2291_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2295
         assign bnn_Add_4Sx2S_4S_1_2295_out1 = bnn_Add_3Sx3S_4S_1_2275_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_2274_out1[1]}}, bnn_N_Mux_2_2_3_1_2274_out1};

         assign bnn_N_Mux_2_2_3_4_2297_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[3], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_1_2270_out1 or bnn_N_Mux_2_2_3_4_2297_in3)
          begin :bnn_N_Mux_2_2_3_4_2297
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2297_out1 = bnn_Minus_2S_2S_1_2270_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2297_out1 = bnn_N_Mux_2_2_3_4_2297_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2298
         assign bnn_Add_3Sx3S_4S_1_2298_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2278_out1[1]}}, bnn_N_Mux_2_2_3_4_2278_out1} + {bnn_Add_2Sx2S_3S_1_2277_out1[2], bnn_Add_2Sx2S_3S_1_2277_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2300
         assign bnn_Add_2Sx2S_3S_1_2300_out1 = {bnn_N_Mux_2_2_3_1_2280_out1[1], bnn_N_Mux_2_2_3_1_2280_out1} + {bnn_N_Mux_2_2_3_1_2279_out1[1], bnn_N_Mux_2_2_3_1_2279_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1815_out1 or bnn_Minus_2S_2S_1_2281_out1)
          begin :bnn_N_Mux_2_2_3_4_2301
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2301_out1 = bnn_Minus_2S_2S_1_2281_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2301_out1 = bnn_N_Mux_2_2_3_1_1815_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1815_out1 or bnn_Minus_2S_2S_1_2281_out1)
          begin :bnn_N_Mux_2_2_3_1_2302
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2302_out1 = bnn_Minus_2S_2S_1_2281_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2302_out1 = bnn_N_Mux_2_2_3_1_1815_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1810_out1 or bnn_Minus_2S_2S_1_2261_out1)
          begin :bnn_N_Mux_2_2_3_1_2303
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2303_out1 = bnn_Minus_2S_2S_1_2261_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2303_out1 = bnn_N_Mux_2_2_3_1_1810_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2304
         assign bnn_Minus_2S_2S_1_2304_out1 = -bnn_N_Mux_2_2_3_1_1820_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1828_out1 or bnn_Minus_2S_2S_4_2267_out1)
          begin :bnn_N_Mux_2_2_3_4_2308
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2308_out1 = bnn_Minus_2S_2S_4_2267_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2308_out1 = bnn_N_Mux_2_2_3_1_1828_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2309
         assign bnn_Add_4Sx2S_5S_1_2309_out1 = {bnn_Add_4Sx2S_4S_1_2286_out1[3], bnn_Add_4Sx2S_4S_1_2286_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2285_out1[1]}}, bnn_N_Mux_2_2_3_4_2285_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2310
         assign bnn_Minus_2S_2S_4_2310_out1 = -bnn_N_Mux_2_2_3_1_1854_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1843_out1 or bnn_Minus_2S_2S_4_2287_out1)
          begin :bnn_N_Mux_2_2_3_4_2311
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2311_out1 = bnn_Minus_2S_2S_4_2287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2311_out1 = bnn_N_Mux_2_2_3_1_1843_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_4Sx2S_5S_1_2289_out1 or bnn_Mod_6Ux32U_7U_4_4991_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2312_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2312_in2 = bnn_Mod_6Ux32U_7U_4_4991_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2312_in2 = {bnn_Add_4Sx2S_5S_1_2289_out1[4], bnn_Add_4Sx2S_5S_1_2289_out1};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_874[6:1] or bnn_N_Mux_2_2_3_4_2288_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2312_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2312_in1 = s_reg_874[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2312_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2288_out1[1]}}, bnn_N_Mux_2_2_3_4_2288_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2312
         assign bnn_Add_6Ux6U_6U_1_2312_out1 = bnn_Add_6Ux6U_6U_1_2312_in2 + bnn_Add_6Ux6U_6U_1_2312_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1843_out1 or bnn_Minus_2S_2S_4_2287_out1)
          begin :bnn_N_Mux_2_2_3_4_2314
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2314_out1 = bnn_Minus_2S_2S_4_2287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2314_out1 = bnn_N_Mux_2_2_3_1_1843_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2315
         assign bnn_Add_4Sx2S_5S_1_2315_out1 = {bnn_Add_4Sx2S_4S_1_2292_out1[3], bnn_Add_4Sx2S_4S_1_2292_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_2291_out1[1]}}, bnn_N_Mux_2_2_3_1_2291_out1};

         // resource: mux_2bx2i
         always @(s_reg_983 or bnn_N_Mux_64_2_2_1_1636_out1[4] or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_2317_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_2317_in3 = s_reg_983;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2317_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[4], 1'b1};
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_939 or bnn_Minus_2S_2S_1_2293_out1 or bnn_N_Mux_2_2_3_1_2317_in3)
          begin :bnn_N_Mux_2_2_3_1_2317
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_1_2317_out1 = bnn_Minus_2S_2S_1_2293_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2317_out1 = bnn_N_Mux_2_2_3_1_2317_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2318
         assign bnn_Add_4Sx2S_4S_1_2318_out1 = bnn_Add_4Sx2S_4S_1_2295_out1 + {{ 2 {bnn_N_Mux_2_2_3_1_2294_out1[1]}}, bnn_N_Mux_2_2_3_1_2294_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2319
         assign bnn_Minus_2S_2S_4_2319_out1 = -bnn_N_Mux_2_4_8_1_1885_in3;

         assign bnn_N_Mux_2_2_3_4_2320_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[4], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_1_2293_out1 or bnn_N_Mux_2_2_3_4_2320_in3)
          begin :bnn_N_Mux_2_2_3_4_2320
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2320_out1 = bnn_Minus_2S_2S_1_2293_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2320_out1 = bnn_N_Mux_2_2_3_4_2320_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2321
         assign bnn_Add_4Sx2S_4S_1_2321_out1 = bnn_Add_3Sx3S_4S_1_2298_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2297_out1[1]}}, bnn_N_Mux_2_2_3_4_2297_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_1_2293_out1 or bnn_N_Mux_2_2_3_4_2320_in3)
          begin :bnn_N_Mux_2_2_3_4_2323
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2323_out1 = bnn_Minus_2S_2S_1_2293_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2323_out1 = bnn_N_Mux_2_2_3_4_2320_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2324
         assign bnn_Add_3Sx3S_4S_1_2324_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2301_out1[1]}}, bnn_N_Mux_2_2_3_4_2301_out1} + {bnn_Add_2Sx2S_3S_1_2300_out1[2], bnn_Add_2Sx2S_3S_1_2300_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2326
         assign bnn_Add_2Sx2S_3S_1_2326_out1 = {bnn_N_Mux_2_2_3_1_2303_out1[1], bnn_N_Mux_2_2_3_1_2303_out1} + {bnn_N_Mux_2_2_3_1_2302_out1[1], bnn_N_Mux_2_2_3_1_2302_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1820_out1 or bnn_Minus_2S_2S_1_2304_out1)
          begin :bnn_N_Mux_2_2_3_4_2327
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2327_out1 = bnn_Minus_2S_2S_1_2304_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2327_out1 = bnn_N_Mux_2_2_3_1_1820_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1820_out1 or bnn_Minus_2S_2S_1_2304_out1)
          begin :bnn_N_Mux_2_2_3_1_2328
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2328_out1 = bnn_Minus_2S_2S_1_2304_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2328_out1 = bnn_N_Mux_2_2_3_1_1820_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1815_out1 or bnn_Minus_2S_2S_1_2281_out1)
          begin :bnn_N_Mux_2_2_3_1_2329
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2329_out1 = bnn_Minus_2S_2S_1_2281_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2329_out1 = bnn_N_Mux_2_2_3_1_1815_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2330
         assign bnn_Minus_2S_2S_1_2330_out1 = -bnn_N_Mux_2_2_3_1_2152_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2331
         assign bnn_Minus_2S_2S_1_2331_out1 = -bnn_N_Mux_2_2_3_1_1825_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2332
         assign bnn_Minus_2S_2S_1_2332_out1 = -bnn_N_Mux_2_2_3_1_1918_out1;

         assign bnn_N_Mux_3_2_6_4_2333_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[7], bnn_N_Mux_64_2_2_1_1636_out1[7]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_2333_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_2333
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_2333_out1_slice = bnn_N_Mux_3_2_6_4_2333_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_2333_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1843_out1 or bnn_Minus_2S_2S_4_2287_out1)
          begin :bnn_N_Mux_2_2_3_4_2334
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2334_out1 = bnn_Minus_2S_2S_4_2287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2334_out1 = bnn_N_Mux_2_2_3_1_1843_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2335
         assign bnn_Add_5Sx4S_6S_1_2335_out1 = {bnn_Add_4Sx2S_5S_1_2309_out1[4], bnn_Add_4Sx2S_5S_1_2309_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2308_out1[1]}}, bnn_N_Mux_2_2_3_4_2308_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1854_out1 or bnn_Minus_2S_2S_4_2310_out1)
          begin :bnn_N_Mux_2_2_3_4_2336
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2336_out1 = bnn_Minus_2S_2S_4_2310_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2336_out1 = bnn_N_Mux_2_2_3_1_1854_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_6Ux6U_6U_1_2312_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4586_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2337_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2337_in2 = bnn_Mod_5Ux32U_7U_1_4586_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2337_in2 = {bnn_Add_6Ux6U_6U_1_2312_out1[4], bnn_Add_6Ux6U_6U_1_2312_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2311_out1 or bnn_LeftShift_9Ux3U_7U_4_4585_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2337_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2337_in1 = bnn_LeftShift_9Ux3U_7U_4_4585_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2337_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2311_out1[1]}}, bnn_N_Mux_2_2_3_4_2311_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2337
         assign bnn_Add_6Ux6U_6U_1_2337_out1 = bnn_Add_6Ux6U_6U_1_2337_in2 + bnn_Add_6Ux6U_6U_1_2337_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2338
         assign bnn_Minus_2S_2S_4_2338_out1 = -bnn_N_Mux_2_2_3_1_1865_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1854_out1 or bnn_Minus_2S_2S_4_2310_out1)
          begin :bnn_N_Mux_2_2_3_4_2339
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2339_out1 = bnn_Minus_2S_2S_4_2310_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2339_out1 = bnn_N_Mux_2_2_3_1_1854_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2340
         assign bnn_Add_5Sx4S_6S_1_2340_out1 = {bnn_Add_4Sx2S_5S_1_2315_out1[4], bnn_Add_4Sx2S_5S_1_2315_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2314_out1[1]}}, bnn_N_Mux_2_2_3_4_2314_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1854_out1 or bnn_Minus_2S_2S_4_2310_out1)
          begin :bnn_N_Mux_2_2_3_4_2342
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2342_out1 = bnn_Minus_2S_2S_4_2310_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2342_out1 = bnn_N_Mux_2_2_3_1_1854_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2343
         assign bnn_Add_4Sx2S_5S_1_2343_out1 = {bnn_Add_4Sx2S_4S_1_2318_out1[3], bnn_Add_4Sx2S_4S_1_2318_out1} + {{ 3 {bnn_N_Mux_2_2_3_1_2317_out1[1]}}, bnn_N_Mux_2_2_3_1_2317_out1};

         assign bnn_N_Mux_2_2_3_4_2345_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[5], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2319_out1 or bnn_N_Mux_2_2_3_4_2345_in3)
          begin :bnn_N_Mux_2_2_3_4_2345
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2345_out1 = bnn_Minus_2S_2S_4_2319_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2345_out1 = bnn_N_Mux_2_2_3_4_2345_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2346
         assign bnn_Add_4Sx2S_4S_1_2346_out1 = bnn_Add_4Sx2S_4S_1_2321_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2320_out1[1]}}, bnn_N_Mux_2_2_3_4_2320_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2347
         assign bnn_Minus_2S_2S_4_2347_out1 = -bnn_N_Mux_2_4_8_1_1896_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2319_out1 or bnn_N_Mux_2_2_3_4_2345_in3)
          begin :bnn_N_Mux_2_2_3_4_2348
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2348_out1 = bnn_Minus_2S_2S_4_2319_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2348_out1 = bnn_N_Mux_2_2_3_4_2345_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2349
         assign bnn_Add_4Sx2S_4S_1_2349_out1 = bnn_Add_3Sx3S_4S_1_2324_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2323_out1[1]}}, bnn_N_Mux_2_2_3_4_2323_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2319_out1 or bnn_N_Mux_2_2_3_4_2345_in3)
          begin :bnn_N_Mux_2_2_3_4_2351
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2351_out1 = bnn_Minus_2S_2S_4_2319_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2351_out1 = bnn_N_Mux_2_2_3_4_2345_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2352
         assign bnn_Add_3Sx3S_4S_1_2352_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2327_out1[1]}}, bnn_N_Mux_2_2_3_4_2327_out1} + {bnn_Add_2Sx2S_3S_1_2326_out1[2], bnn_Add_2Sx2S_3S_1_2326_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2354
         assign bnn_Add_2Sx2S_3S_1_2354_out1 = {bnn_N_Mux_2_2_3_1_2329_out1[1], bnn_N_Mux_2_2_3_1_2329_out1} + {bnn_N_Mux_2_2_3_1_2328_out1[1], bnn_N_Mux_2_2_3_1_2328_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2152_out1 or bnn_Minus_2S_2S_1_2330_out1)
          begin :bnn_N_Mux_2_2_3_4_2355
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2355_out1 = bnn_Minus_2S_2S_1_2330_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2355_out1 = bnn_N_Mux_2_2_3_1_2152_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_Minus_2S_2S_1_2331_out1)
          begin :bnn_N_Mux_2_2_3_4_2356
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2356_out1 = bnn_Minus_2S_2S_1_2331_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2356_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1918_out1 or bnn_Minus_2S_2S_1_2332_out1)
          begin :bnn_N_Mux_2_2_3_4_2357
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2357_out1 = bnn_Minus_2S_2S_1_2332_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2357_out1 = bnn_N_Mux_2_2_3_1_1918_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2358
         assign bnn_Minus_2S_2S_1_2358_out1 = -bnn_N_Mux_2_2_3_1_1840_out1;

         assign bnn_N_Mux_3_2_6_4_2361_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[8], bnn_N_Mux_64_2_2_1_1636_out1[8]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_2361_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_2361
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_2361_out1_slice = bnn_N_Mux_3_2_6_4_2361_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_2361_out1_slice = 2'd0;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2335_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4595_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2362_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2362_in2 = bnn_Mod_5Ux32U_7U_1_4595_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2362_in2 = {bnn_Add_5Sx4S_6S_1_2335_out1[4], bnn_Add_5Sx4S_6S_1_2335_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2334_out1 or bnn_LeftShift_9Ux3U_7U_4_4594_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2362_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2362_in1 = bnn_LeftShift_9Ux3U_7U_4_4594_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2362_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2334_out1[1]}}, bnn_N_Mux_2_2_3_4_2334_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2362
         assign bnn_Add_6Ux6U_6U_1_2362_out1 = bnn_Add_6Ux6U_6U_1_2362_in2 + bnn_Add_6Ux6U_6U_1_2362_in1;

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2363
         assign bnn_Add_5Sx4S_6S_1_2363_out1 = {bnn_Add_6Ux6U_6U_1_2337_out1[4], bnn_Add_6Ux6U_6U_1_2337_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2336_out1[1]}}, bnn_N_Mux_2_2_3_4_2336_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1865_out1 or bnn_Minus_2S_2S_4_2338_out1)
          begin :bnn_N_Mux_2_2_3_4_2364
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2364_out1 = bnn_Minus_2S_2S_4_2338_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2364_out1 = bnn_N_Mux_2_2_3_1_1865_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2340_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4604_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2365_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2365_in2 = bnn_Mod_5Ux32U_7U_1_4604_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2365_in2 = {bnn_Add_5Sx4S_6S_1_2340_out1[4], bnn_Add_5Sx4S_6S_1_2340_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2339_out1 or bnn_LeftShift_9Ux3U_7U_4_4603_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2365_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2365_in1 = bnn_LeftShift_9Ux3U_7U_4_4603_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2365_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2339_out1[1]}}, bnn_N_Mux_2_2_3_4_2339_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2365
         assign bnn_Add_6Ux6U_6U_1_2365_out1 = bnn_Add_6Ux6U_6U_1_2365_in2 + bnn_Add_6Ux6U_6U_1_2365_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2366
         assign bnn_Minus_2S_2S_4_2366_out1 = -bnn_N_Mux_2_2_3_1_1876_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1865_out1 or bnn_Minus_2S_2S_4_2338_out1)
          begin :bnn_N_Mux_2_2_3_4_2367
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2367_out1 = bnn_Minus_2S_2S_4_2338_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2367_out1 = bnn_N_Mux_2_2_3_1_1865_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2368
         assign bnn_Add_5Sx4S_6S_1_2368_out1 = {bnn_Add_4Sx2S_5S_1_2343_out1[4], bnn_Add_4Sx2S_5S_1_2343_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2342_out1[1]}}, bnn_N_Mux_2_2_3_4_2342_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1865_out1 or bnn_Minus_2S_2S_4_2338_out1)
          begin :bnn_N_Mux_2_2_3_4_2370
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2370_out1 = bnn_Minus_2S_2S_4_2338_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2370_out1 = bnn_N_Mux_2_2_3_1_1865_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2371
         assign bnn_Add_4Sx2S_5S_1_2371_out1 = {bnn_Add_4Sx2S_4S_1_2346_out1[3], bnn_Add_4Sx2S_4S_1_2346_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2345_out1[1]}}, bnn_N_Mux_2_2_3_4_2345_out1};

         assign bnn_N_Mux_2_2_3_4_2373_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[6], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2347_out1 or bnn_N_Mux_2_2_3_4_2373_in3)
          begin :bnn_N_Mux_2_2_3_4_2373
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2373_out1 = bnn_Minus_2S_2S_4_2347_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2373_out1 = bnn_N_Mux_2_2_3_4_2373_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2374
         assign bnn_Add_4Sx2S_4S_1_2374_out1 = bnn_Add_4Sx2S_4S_1_2349_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2348_out1[1]}}, bnn_N_Mux_2_2_3_4_2348_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2375
         assign bnn_Minus_2S_2S_4_2375_out1 = -bnn_N_Mux_2_4_8_1_1907_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2347_out1 or bnn_N_Mux_2_2_3_4_2373_in3)
          begin :bnn_N_Mux_2_2_3_4_2376
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2376_out1 = bnn_Minus_2S_2S_4_2347_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2376_out1 = bnn_N_Mux_2_2_3_4_2373_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2377
         assign bnn_Add_4Sx2S_4S_1_2377_out1 = bnn_Add_3Sx3S_4S_1_2352_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2351_out1[1]}}, bnn_N_Mux_2_2_3_4_2351_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2347_out1 or bnn_N_Mux_2_2_3_4_2373_in3)
          begin :bnn_N_Mux_2_2_3_4_2379
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2379_out1 = bnn_Minus_2S_2S_4_2347_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2379_out1 = bnn_N_Mux_2_2_3_4_2373_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2380
         assign bnn_Add_3Sx3S_4S_1_2380_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2355_out1[1]}}, bnn_N_Mux_2_2_3_4_2355_out1} + {bnn_Add_2Sx2S_3S_1_2354_out1[2], bnn_Add_2Sx2S_3S_1_2354_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2381
         assign bnn_Minus_2S_2S_4_2381_out1 = -bnn_N_Mux_3_2_6_4_2333_out1_slice;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2382
         assign bnn_Add_2Sx2S_3S_1_2382_out1 = {bnn_N_Mux_2_2_3_4_2357_out1[1], bnn_N_Mux_2_2_3_4_2357_out1} + {bnn_N_Mux_2_2_3_4_2356_out1[1], bnn_N_Mux_2_2_3_4_2356_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_Minus_2S_2S_1_2358_out1)
          begin :bnn_N_Mux_2_2_3_4_2383
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2383_out1 = bnn_Minus_2S_2S_1_2358_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2383_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_Minus_2S_2S_1_2358_out1)
          begin :bnn_N_Mux_2_2_3_1_2384
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2384_out1 = bnn_Minus_2S_2S_1_2358_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2384_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1825_out1 or bnn_Minus_2S_2S_1_2331_out1)
          begin :bnn_N_Mux_2_2_3_1_2385
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2385_out1 = bnn_Minus_2S_2S_1_2331_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2385_out1 = bnn_N_Mux_2_2_3_1_1825_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2386
         assign bnn_Minus_2S_2S_1_2386_out1 = -bnn_N_Mux_2_2_3_1_1851_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_0_if_1_dout_wire or bnn_Mul_30Sx12S_30S_1_191_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2389_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2389_in2 = {bnn_Mul_30Sx12S_30S_1_191_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2389_in2 = {{ 5 {fixed_buffer_0_if_1_dout_wire[11]}}, fixed_buffer_0_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_2362_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2389_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2389_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2389_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_2362_out1[4]}}, bnn_Add_6Ux6U_6U_1_2362_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2389
         assign bnn_Add_17Sx16S_17S_1_2389_out1 = bnn_Add_17Sx16S_17S_1_2389_in2 + {bnn_Add_17Sx16S_17S_1_2389_in1[15], bnn_Add_17Sx16S_17S_1_2389_in1};

         // resource: mux_17bx2i
         always @(fixed_buffer_1_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4715_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2390_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2390_in2 = {bnn_Mul_16Sx12S_19S_4_4715_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2390_in2 = {{ 5 {fixed_buffer_1_if_1_dout_wire[11]}}, fixed_buffer_1_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2363_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2390_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2390_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2390_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2363_out1[4]}}, bnn_Add_5Sx4S_6S_1_2363_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2390
         assign bnn_Add_17Sx16S_17S_1_2390_out1 = bnn_Add_17Sx16S_17S_1_2390_in2 + {bnn_Add_17Sx16S_17S_1_2390_in1[15], bnn_Add_17Sx16S_17S_1_2390_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2391
         assign bnn_Add_5Sx4S_6S_1_2391_out1 = {bnn_Add_6Ux6U_6U_1_2365_out1[4], bnn_Add_6Ux6U_6U_1_2365_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2364_out1[1]}}, bnn_N_Mux_2_2_3_4_2364_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1876_out1 or bnn_Minus_2S_2S_4_2366_out1)
          begin :bnn_N_Mux_2_2_3_4_2392
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2392_out1 = bnn_Minus_2S_2S_4_2366_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2392_out1 = bnn_N_Mux_2_2_3_1_1876_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2368_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4613_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2393_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2393_in2 = bnn_Mod_5Ux32U_7U_1_4613_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2393_in2 = {bnn_Add_5Sx4S_6S_1_2368_out1[4], bnn_Add_5Sx4S_6S_1_2368_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2367_out1 or bnn_LeftShift_9Ux3U_7U_4_4612_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2393_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2393_in1 = bnn_LeftShift_9Ux3U_7U_4_4612_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2393_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2367_out1[1]}}, bnn_N_Mux_2_2_3_4_2367_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2393
         assign bnn_Add_6Ux6U_6U_1_2393_out1 = bnn_Add_6Ux6U_6U_1_2393_in2 + bnn_Add_6Ux6U_6U_1_2393_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2394
         assign bnn_Minus_2S_2S_4_2394_out1 = -bnn_N_Mux_2_2_3_1_1887_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1876_out1 or bnn_Minus_2S_2S_4_2366_out1)
          begin :bnn_N_Mux_2_2_3_4_2395
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2395_out1 = bnn_Minus_2S_2S_4_2366_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2395_out1 = bnn_N_Mux_2_2_3_1_1876_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2396
         assign bnn_Add_5Sx4S_6S_1_2396_out1 = {bnn_Add_4Sx2S_5S_1_2371_out1[4], bnn_Add_4Sx2S_5S_1_2371_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2370_out1[1]}}, bnn_N_Mux_2_2_3_4_2370_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1876_out1 or bnn_Minus_2S_2S_4_2366_out1)
          begin :bnn_N_Mux_2_2_3_4_2398
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2398_out1 = bnn_Minus_2S_2S_4_2366_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2398_out1 = bnn_N_Mux_2_2_3_1_1876_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2399
         assign bnn_Add_4Sx2S_5S_1_2399_out1 = {bnn_Add_4Sx2S_4S_1_2374_out1[3], bnn_Add_4Sx2S_4S_1_2374_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2373_out1[1]}}, bnn_N_Mux_2_2_3_4_2373_out1};

         assign bnn_N_Mux_2_2_3_4_2401_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[7], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2375_out1 or bnn_N_Mux_2_2_3_4_2401_in3)
          begin :bnn_N_Mux_2_2_3_4_2401
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2401_out1 = bnn_Minus_2S_2S_4_2375_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2401_out1 = bnn_N_Mux_2_2_3_4_2401_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2402
         assign bnn_Add_4Sx2S_4S_1_2402_out1 = bnn_Add_4Sx2S_4S_1_2377_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2376_out1[1]}}, bnn_N_Mux_2_2_3_4_2376_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2403
         assign bnn_Minus_2S_2S_4_2403_out1 = -bnn_N_Mux_3_2_6_4_2361_out1_slice;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2375_out1 or bnn_N_Mux_2_2_3_4_2401_in3)
          begin :bnn_N_Mux_2_2_3_4_2404
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2404_out1 = bnn_Minus_2S_2S_4_2375_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2404_out1 = bnn_N_Mux_2_2_3_4_2401_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2405
         assign bnn_Add_4Sx2S_4S_1_2405_out1 = bnn_Add_3Sx3S_4S_1_2380_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2379_out1[1]}}, bnn_N_Mux_2_2_3_4_2379_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2406
         assign bnn_Minus_2S_2S_4_2406_out1 = -bnn_N_Mux_2_4_8_1_1928_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2381_out1 or bnn_N_Mux_3_2_6_4_2333_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2407
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2407_out1 = bnn_Minus_2S_2S_4_2381_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2407_out1 = bnn_N_Mux_3_2_6_4_2333_out1_slice;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2408
         assign bnn_Add_3Sx3S_4S_1_2408_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2383_out1[1]}}, bnn_N_Mux_2_2_3_4_2383_out1} + {bnn_Add_2Sx2S_3S_1_2382_out1[2], bnn_Add_2Sx2S_3S_1_2382_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2410
         assign bnn_Add_2Sx2S_3S_1_2410_out1 = {bnn_N_Mux_2_2_3_1_2385_out1[1], bnn_N_Mux_2_2_3_1_2385_out1} + {bnn_N_Mux_2_2_3_1_2384_out1[1], bnn_N_Mux_2_2_3_1_2384_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_Minus_2S_2S_1_2386_out1)
          begin :bnn_N_Mux_2_2_3_4_2411
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2411_out1 = bnn_Minus_2S_2S_1_2386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2411_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_Minus_2S_2S_1_2386_out1)
          begin :bnn_N_Mux_2_2_3_1_2412
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2412_out1 = bnn_Minus_2S_2S_1_2386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2412_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1840_out1 or bnn_Minus_2S_2S_1_2358_out1)
          begin :bnn_N_Mux_2_2_3_1_2413
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2413_out1 = bnn_Minus_2S_2S_1_2358_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2413_out1 = bnn_N_Mux_2_2_3_1_1840_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2414
         assign bnn_Minus_2S_2S_1_2414_out1 = -bnn_N_Mux_2_2_3_1_1862_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_2_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4724_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2417_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2417_in2 = {bnn_Mul_16Sx12S_19S_4_4724_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2417_in2 = {{ 5 {fixed_buffer_2_if_1_dout_wire[11]}}, fixed_buffer_2_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2391_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2417_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2417_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2417_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2391_out1[4]}}, bnn_Add_5Sx4S_6S_1_2391_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2417
         assign bnn_Add_17Sx16S_17S_1_2417_out1 = bnn_Add_17Sx16S_17S_1_2417_in2 + {bnn_Add_17Sx16S_17S_1_2417_in1[15], bnn_Add_17Sx16S_17S_1_2417_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2418
         assign bnn_Add_5Sx4S_6S_1_2418_out1 = {bnn_Add_6Ux6U_6U_1_2393_out1[4], bnn_Add_6Ux6U_6U_1_2393_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2392_out1[1]}}, bnn_N_Mux_2_2_3_4_2392_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1887_out1 or bnn_Minus_2S_2S_4_2394_out1)
          begin :bnn_N_Mux_2_2_3_4_2419
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2419_out1 = bnn_Minus_2S_2S_4_2394_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2419_out1 = bnn_N_Mux_2_2_3_1_1887_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2396_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4622_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2420_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2420_in2 = bnn_Mod_5Ux32U_7U_1_4622_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2420_in2 = {bnn_Add_5Sx4S_6S_1_2396_out1[4], bnn_Add_5Sx4S_6S_1_2396_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2395_out1 or bnn_LeftShift_9Ux3U_7U_4_4621_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2420_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2420_in1 = bnn_LeftShift_9Ux3U_7U_4_4621_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2420_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2395_out1[1]}}, bnn_N_Mux_2_2_3_4_2395_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2420
         assign bnn_Add_6Ux6U_6U_1_2420_out1 = bnn_Add_6Ux6U_6U_1_2420_in2 + bnn_Add_6Ux6U_6U_1_2420_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2421
         assign bnn_Minus_2S_2S_4_2421_out1 = -bnn_N_Mux_2_2_3_1_1898_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1887_out1 or bnn_Minus_2S_2S_4_2394_out1)
          begin :bnn_N_Mux_2_2_3_4_2422
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2422_out1 = bnn_Minus_2S_2S_4_2394_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2422_out1 = bnn_N_Mux_2_2_3_1_1887_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2423
         assign bnn_Add_5Sx4S_6S_1_2423_out1 = {bnn_Add_4Sx2S_5S_1_2399_out1[4], bnn_Add_4Sx2S_5S_1_2399_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2398_out1[1]}}, bnn_N_Mux_2_2_3_4_2398_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1887_out1 or bnn_Minus_2S_2S_4_2394_out1)
          begin :bnn_N_Mux_2_2_3_4_2425
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2425_out1 = bnn_Minus_2S_2S_4_2394_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2425_out1 = bnn_N_Mux_2_2_3_1_1887_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2426
         assign bnn_Add_4Sx2S_5S_1_2426_out1 = {bnn_Add_4Sx2S_4S_1_2402_out1[3], bnn_Add_4Sx2S_4S_1_2402_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2401_out1[1]}}, bnn_N_Mux_2_2_3_4_2401_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2403_out1 or bnn_N_Mux_3_2_6_4_2361_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2428
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2428_out1 = bnn_Minus_2S_2S_4_2403_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2428_out1 = bnn_N_Mux_3_2_6_4_2361_out1_slice;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2429
         assign bnn_Add_4Sx2S_4S_1_2429_out1 = bnn_Add_4Sx2S_4S_1_2405_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2404_out1[1]}}, bnn_N_Mux_2_2_3_4_2404_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2430
         assign bnn_Minus_2S_2S_4_2430_out1 = -bnn_N_Mux_2_4_8_1_1939_in3;

         assign bnn_N_Mux_2_2_3_4_2431_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[8], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2406_out1 or bnn_N_Mux_2_2_3_4_2431_in3)
          begin :bnn_N_Mux_2_2_3_4_2431
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2431_out1 = bnn_Minus_2S_2S_4_2406_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2431_out1 = bnn_N_Mux_2_2_3_4_2431_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2432
         assign bnn_Add_4Sx3S_4S_1_2432_out1 = bnn_Add_3Sx3S_4S_1_2408_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2407_out1[1]}}, bnn_N_Mux_2_2_3_4_2407_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2406_out1 or bnn_N_Mux_2_2_3_4_2431_in3)
          begin :bnn_N_Mux_2_2_3_4_2434
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2434_out1 = bnn_Minus_2S_2S_4_2406_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2434_out1 = bnn_N_Mux_2_2_3_4_2431_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2435
         assign bnn_Add_3Sx3S_4S_1_2435_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2411_out1[1]}}, bnn_N_Mux_2_2_3_4_2411_out1} + {bnn_Add_2Sx2S_3S_1_2410_out1[2], bnn_Add_2Sx2S_3S_1_2410_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2437
         assign bnn_Add_2Sx2S_3S_1_2437_out1 = {bnn_N_Mux_2_2_3_1_2413_out1[1], bnn_N_Mux_2_2_3_1_2413_out1} + {bnn_N_Mux_2_2_3_1_2412_out1[1], bnn_N_Mux_2_2_3_1_2412_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_Minus_2S_2S_1_2414_out1)
          begin :bnn_N_Mux_2_2_3_4_2438
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2438_out1 = bnn_Minus_2S_2S_1_2414_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2438_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_Minus_2S_2S_1_2414_out1)
          begin :bnn_N_Mux_2_2_3_1_2439
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2439_out1 = bnn_Minus_2S_2S_1_2414_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2439_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1851_out1 or bnn_Minus_2S_2S_1_2386_out1)
          begin :bnn_N_Mux_2_2_3_1_2440
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2440_out1 = bnn_Minus_2S_2S_1_2386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2440_out1 = bnn_N_Mux_2_2_3_1_1851_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2441
         assign bnn_Minus_2S_2S_1_2441_out1 = -bnn_N_Mux_2_2_3_1_1873_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_3_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4732_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2444_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2444_in2 = {bnn_Mul_16Sx12S_19S_4_4732_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2444_in2 = {{ 5 {fixed_buffer_3_if_1_dout_wire[11]}}, fixed_buffer_3_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2418_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2444_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2444_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2444_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2418_out1[4]}}, bnn_Add_5Sx4S_6S_1_2418_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2444
         assign bnn_Add_17Sx16S_17S_1_2444_out1 = bnn_Add_17Sx16S_17S_1_2444_in2 + {bnn_Add_17Sx16S_17S_1_2444_in1[15], bnn_Add_17Sx16S_17S_1_2444_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2445
         assign bnn_Add_5Sx4S_6S_1_2445_out1 = {bnn_Add_6Ux6U_6U_1_2420_out1[4], bnn_Add_6Ux6U_6U_1_2420_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2419_out1[1]}}, bnn_N_Mux_2_2_3_4_2419_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1898_out1 or bnn_Minus_2S_2S_4_2421_out1)
          begin :bnn_N_Mux_2_2_3_4_2446
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2446_out1 = bnn_Minus_2S_2S_4_2421_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2446_out1 = bnn_N_Mux_2_2_3_1_1898_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2423_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4631_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2447_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2447_in2 = bnn_Mod_5Ux32U_7U_1_4631_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2447_in2 = {bnn_Add_5Sx4S_6S_1_2423_out1[4], bnn_Add_5Sx4S_6S_1_2423_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2422_out1 or bnn_LeftShift_9Ux3U_7U_4_4630_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2447_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2447_in1 = bnn_LeftShift_9Ux3U_7U_4_4630_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2447_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2422_out1[1]}}, bnn_N_Mux_2_2_3_4_2422_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2447
         assign bnn_Add_6Ux6U_6U_1_2447_out1 = bnn_Add_6Ux6U_6U_1_2447_in2 + bnn_Add_6Ux6U_6U_1_2447_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2448
         assign bnn_Minus_2S_2S_4_2448_out1 = -bnn_N_Mux_2_2_3_1_1909_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1898_out1 or bnn_Minus_2S_2S_4_2421_out1)
          begin :bnn_N_Mux_2_2_3_4_2449
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2449_out1 = bnn_Minus_2S_2S_4_2421_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2449_out1 = bnn_N_Mux_2_2_3_1_1898_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2450
         assign bnn_Add_5Sx4S_6S_1_2450_out1 = {bnn_Add_4Sx2S_5S_1_2426_out1[4], bnn_Add_4Sx2S_5S_1_2426_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2425_out1[1]}}, bnn_N_Mux_2_2_3_4_2425_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1898_out1 or bnn_Minus_2S_2S_4_2421_out1)
          begin :bnn_N_Mux_2_2_3_4_2452
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2452_out1 = bnn_Minus_2S_2S_4_2421_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2452_out1 = bnn_N_Mux_2_2_3_1_1898_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2453
         assign bnn_Add_4Sx2S_5S_1_2453_out1 = {bnn_Add_4Sx2S_4S_1_2429_out1[3], bnn_Add_4Sx2S_4S_1_2429_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2428_out1[1]}}, bnn_N_Mux_2_2_3_4_2428_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2454
         assign bnn_Minus_2S_2S_4_2454_out1 = -bnn_N_Mux_2_2_3_1_2173_out1;

         assign bnn_N_Mux_2_2_3_4_2455_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[9], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2430_out1 or bnn_N_Mux_2_2_3_4_2455_in3)
          begin :bnn_N_Mux_2_2_3_4_2455
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2455_out1 = bnn_Minus_2S_2S_4_2430_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2455_out1 = bnn_N_Mux_2_2_3_4_2455_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2456
         assign bnn_Add_4Sx3S_4S_1_2456_out1 = bnn_Add_4Sx3S_4S_1_2432_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2431_out1[1]}}, bnn_N_Mux_2_2_3_4_2431_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2457
         assign bnn_Minus_2S_2S_4_2457_out1 = -bnn_N_Mux_2_4_8_1_1950_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2430_out1 or bnn_N_Mux_2_2_3_4_2455_in3)
          begin :bnn_N_Mux_2_2_3_4_2458
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2458_out1 = bnn_Minus_2S_2S_4_2430_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2458_out1 = bnn_N_Mux_2_2_3_4_2455_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2459
         assign bnn_Add_4Sx2S_4S_1_2459_out1 = bnn_Add_3Sx3S_4S_1_2435_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2434_out1[1]}}, bnn_N_Mux_2_2_3_4_2434_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2430_out1 or bnn_N_Mux_2_2_3_4_2455_in3)
          begin :bnn_N_Mux_2_2_3_4_2461
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2461_out1 = bnn_Minus_2S_2S_4_2430_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2461_out1 = bnn_N_Mux_2_2_3_4_2455_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2462
         assign bnn_Add_3Sx3S_4S_1_2462_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2438_out1[1]}}, bnn_N_Mux_2_2_3_4_2438_out1} + {bnn_Add_2Sx2S_3S_1_2437_out1[2], bnn_Add_2Sx2S_3S_1_2437_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2464
         assign bnn_Add_2Sx2S_3S_1_2464_out1 = {bnn_N_Mux_2_2_3_1_2440_out1[1], bnn_N_Mux_2_2_3_1_2440_out1} + {bnn_N_Mux_2_2_3_1_2439_out1[1], bnn_N_Mux_2_2_3_1_2439_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_Minus_2S_2S_1_2441_out1)
          begin :bnn_N_Mux_2_2_3_4_2465
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2465_out1 = bnn_Minus_2S_2S_1_2441_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2465_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_Minus_2S_2S_1_2441_out1)
          begin :bnn_N_Mux_2_2_3_1_2466
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2466_out1 = bnn_Minus_2S_2S_1_2441_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2466_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1862_out1 or bnn_Minus_2S_2S_1_2414_out1)
          begin :bnn_N_Mux_2_2_3_1_2467
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2467_out1 = bnn_Minus_2S_2S_1_2414_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2467_out1 = bnn_N_Mux_2_2_3_1_1862_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2468
         assign bnn_Minus_2S_2S_1_2468_out1 = -bnn_N_Mux_2_2_3_1_1884_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_4_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4739_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2471_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2471_in2 = {bnn_Mul_16Sx12S_19S_4_4739_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2471_in2 = {{ 5 {fixed_buffer_4_if_1_dout_wire[11]}}, fixed_buffer_4_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2445_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2471_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2471_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2471_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2445_out1[4]}}, bnn_Add_5Sx4S_6S_1_2445_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2471
         assign bnn_Add_17Sx16S_17S_1_2471_out1 = bnn_Add_17Sx16S_17S_1_2471_in2 + {bnn_Add_17Sx16S_17S_1_2471_in1[15], bnn_Add_17Sx16S_17S_1_2471_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2472
         assign bnn_Add_5Sx4S_6S_1_2472_out1 = {bnn_Add_6Ux6U_6U_1_2447_out1[4], bnn_Add_6Ux6U_6U_1_2447_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2446_out1[1]}}, bnn_N_Mux_2_2_3_4_2446_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1909_out1 or bnn_Minus_2S_2S_4_2448_out1)
          begin :bnn_N_Mux_2_2_3_4_2473
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2473_out1 = bnn_Minus_2S_2S_4_2448_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2473_out1 = bnn_N_Mux_2_2_3_1_1909_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2450_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4640_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2474_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2474_in2 = bnn_Mod_5Ux32U_7U_1_4640_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2474_in2 = {bnn_Add_5Sx4S_6S_1_2450_out1[4], bnn_Add_5Sx4S_6S_1_2450_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2449_out1 or bnn_LeftShift_9Ux3U_7U_4_4639_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2474_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2474_in1 = bnn_LeftShift_9Ux3U_7U_4_4639_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2474_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2449_out1[1]}}, bnn_N_Mux_2_2_3_4_2449_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2474
         assign bnn_Add_6Ux6U_6U_1_2474_out1 = bnn_Add_6Ux6U_6U_1_2474_in2 + bnn_Add_6Ux6U_6U_1_2474_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2475
         assign bnn_Minus_2S_2S_4_2475_out1 = -bnn_N_Mux_2_2_3_1_2161_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1909_out1 or bnn_Minus_2S_2S_4_2448_out1)
          begin :bnn_N_Mux_2_2_3_4_2476
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2476_out1 = bnn_Minus_2S_2S_4_2448_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2476_out1 = bnn_N_Mux_2_2_3_1_1909_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2477
         assign bnn_Add_5Sx4S_6S_1_2477_out1 = {bnn_Add_4Sx2S_5S_1_2453_out1[4], bnn_Add_4Sx2S_5S_1_2453_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2452_out1[1]}}, bnn_N_Mux_2_2_3_4_2452_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2478
         assign bnn_Minus_2S_2S_4_2478_out1 = -bnn_N_Mux_2_2_3_1_1930_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2173_out1 or bnn_Minus_2S_2S_4_2454_out1)
          begin :bnn_N_Mux_2_2_3_4_2479
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2479_out1 = bnn_Minus_2S_2S_4_2454_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2479_out1 = bnn_N_Mux_2_2_3_1_2173_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2480
         assign bnn_Add_4Sx2S_5S_1_2480_out1 = {bnn_Add_4Sx3S_4S_1_2456_out1[3], bnn_Add_4Sx3S_4S_1_2456_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2455_out1[1]}}, bnn_N_Mux_2_2_3_4_2455_out1};

         assign bnn_N_Mux_2_2_3_4_2482_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[10], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2457_out1 or bnn_N_Mux_2_2_3_4_2482_in3)
          begin :bnn_N_Mux_2_2_3_4_2482
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2482_out1 = bnn_Minus_2S_2S_4_2457_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2482_out1 = bnn_N_Mux_2_2_3_4_2482_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2483
         assign bnn_Add_4Sx2S_4S_1_2483_out1 = bnn_Add_4Sx2S_4S_1_2459_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2458_out1[1]}}, bnn_N_Mux_2_2_3_4_2458_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2484
         assign bnn_Minus_2S_2S_4_2484_out1 = -bnn_N_Mux_2_4_8_1_1961_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2457_out1 or bnn_N_Mux_2_2_3_4_2482_in3)
          begin :bnn_N_Mux_2_2_3_4_2485
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2485_out1 = bnn_Minus_2S_2S_4_2457_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2485_out1 = bnn_N_Mux_2_2_3_4_2482_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2486
         assign bnn_Add_4Sx2S_4S_1_2486_out1 = bnn_Add_3Sx3S_4S_1_2462_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2461_out1[1]}}, bnn_N_Mux_2_2_3_4_2461_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2457_out1 or bnn_N_Mux_2_2_3_4_2482_in3)
          begin :bnn_N_Mux_2_2_3_4_2488
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2488_out1 = bnn_Minus_2S_2S_4_2457_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2488_out1 = bnn_N_Mux_2_2_3_4_2482_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2489
         assign bnn_Add_3Sx3S_4S_1_2489_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2465_out1[1]}}, bnn_N_Mux_2_2_3_4_2465_out1} + {bnn_Add_2Sx2S_3S_1_2464_out1[2], bnn_Add_2Sx2S_3S_1_2464_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2491
         assign bnn_Add_2Sx2S_3S_1_2491_out1 = {bnn_N_Mux_2_2_3_1_2467_out1[1], bnn_N_Mux_2_2_3_1_2467_out1} + {bnn_N_Mux_2_2_3_1_2466_out1[1], bnn_N_Mux_2_2_3_1_2466_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_Minus_2S_2S_1_2468_out1)
          begin :bnn_N_Mux_2_2_3_4_2492
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2492_out1 = bnn_Minus_2S_2S_1_2468_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2492_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_Minus_2S_2S_1_2468_out1)
          begin :bnn_N_Mux_2_2_3_1_2493
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2493_out1 = bnn_Minus_2S_2S_1_2468_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2493_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1873_out1 or bnn_Minus_2S_2S_1_2441_out1)
          begin :bnn_N_Mux_2_2_3_1_2494
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2494_out1 = bnn_Minus_2S_2S_1_2441_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2494_out1 = bnn_N_Mux_2_2_3_1_1873_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2495
         assign bnn_Minus_2S_2S_1_2495_out1 = -bnn_N_Mux_2_2_3_1_1895_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_5_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4745_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2498_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2498_in2 = {bnn_Mul_16Sx12S_19S_4_4745_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2498_in2 = {{ 5 {fixed_buffer_5_if_1_dout_wire[11]}}, fixed_buffer_5_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2472_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2498_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2498_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2498_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2472_out1[4]}}, bnn_Add_5Sx4S_6S_1_2472_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2498
         assign bnn_Add_17Sx16S_17S_1_2498_out1 = bnn_Add_17Sx16S_17S_1_2498_in2 + {bnn_Add_17Sx16S_17S_1_2498_in1[15], bnn_Add_17Sx16S_17S_1_2498_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2499
         assign bnn_Add_5Sx4S_6S_1_2499_out1 = {bnn_Add_6Ux6U_6U_1_2474_out1[4], bnn_Add_6Ux6U_6U_1_2474_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2473_out1[1]}}, bnn_N_Mux_2_2_3_4_2473_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2161_out1 or bnn_Minus_2S_2S_4_2475_out1)
          begin :bnn_N_Mux_2_2_3_4_2500
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2500_out1 = bnn_Minus_2S_2S_4_2475_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2500_out1 = bnn_N_Mux_2_2_3_1_2161_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2477_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4649_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2501_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2501_in2 = bnn_Mod_5Ux32U_7U_1_4649_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2501_in2 = {bnn_Add_5Sx4S_6S_1_2477_out1[4], bnn_Add_5Sx4S_6S_1_2477_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2476_out1 or bnn_LeftShift_9Ux3U_7U_4_4648_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2501_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2501_in1 = bnn_LeftShift_9Ux3U_7U_4_4648_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2501_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2476_out1[1]}}, bnn_N_Mux_2_2_3_4_2476_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2501
         assign bnn_Add_6Ux6U_6U_1_2501_out1 = bnn_Add_6Ux6U_6U_1_2501_in2 + bnn_Add_6Ux6U_6U_1_2501_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2502
         assign bnn_Minus_2S_2S_4_2502_out1 = -bnn_N_Mux_2_2_3_1_1941_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1930_out1 or bnn_Minus_2S_2S_4_2478_out1)
          begin :bnn_N_Mux_2_2_3_4_2503
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2503_out1 = bnn_Minus_2S_2S_4_2478_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2503_out1 = bnn_N_Mux_2_2_3_1_1930_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2504
         assign bnn_Add_5Sx4S_6S_1_2504_out1 = {bnn_Add_4Sx2S_5S_1_2480_out1[4], bnn_Add_4Sx2S_5S_1_2480_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2479_out1[1]}}, bnn_N_Mux_2_2_3_4_2479_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1930_out1 or bnn_Minus_2S_2S_4_2478_out1)
          begin :bnn_N_Mux_2_2_3_4_2506
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2506_out1 = bnn_Minus_2S_2S_4_2478_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2506_out1 = bnn_N_Mux_2_2_3_1_1930_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2507
         assign bnn_Add_4Sx2S_5S_1_2507_out1 = {bnn_Add_4Sx2S_4S_1_2483_out1[3], bnn_Add_4Sx2S_4S_1_2483_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2482_out1[1]}}, bnn_N_Mux_2_2_3_4_2482_out1};

         assign bnn_N_Mux_2_2_3_4_2509_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[11], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2484_out1 or bnn_N_Mux_2_2_3_4_2509_in3)
          begin :bnn_N_Mux_2_2_3_4_2509
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2509_out1 = bnn_Minus_2S_2S_4_2484_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2509_out1 = bnn_N_Mux_2_2_3_4_2509_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2510
         assign bnn_Add_4Sx2S_4S_1_2510_out1 = bnn_Add_4Sx2S_4S_1_2486_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2485_out1[1]}}, bnn_N_Mux_2_2_3_4_2485_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2511
         assign bnn_Minus_2S_2S_4_2511_out1 = -bnn_N_Mux_2_4_8_1_1972_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2484_out1 or bnn_N_Mux_2_2_3_4_2509_in3)
          begin :bnn_N_Mux_2_2_3_4_2512
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2512_out1 = bnn_Minus_2S_2S_4_2484_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2512_out1 = bnn_N_Mux_2_2_3_4_2509_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2513
         assign bnn_Add_4Sx2S_4S_1_2513_out1 = bnn_Add_3Sx3S_4S_1_2489_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2488_out1[1]}}, bnn_N_Mux_2_2_3_4_2488_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2484_out1 or bnn_N_Mux_2_2_3_4_2509_in3)
          begin :bnn_N_Mux_2_2_3_4_2515
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2515_out1 = bnn_Minus_2S_2S_4_2484_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2515_out1 = bnn_N_Mux_2_2_3_4_2509_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2516
         assign bnn_Add_3Sx3S_4S_1_2516_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2492_out1[1]}}, bnn_N_Mux_2_2_3_4_2492_out1} + {bnn_Add_2Sx2S_3S_1_2491_out1[2], bnn_Add_2Sx2S_3S_1_2491_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2518
         assign bnn_Add_2Sx2S_3S_1_2518_out1 = {bnn_N_Mux_2_2_3_1_2494_out1[1], bnn_N_Mux_2_2_3_1_2494_out1} + {bnn_N_Mux_2_2_3_1_2493_out1[1], bnn_N_Mux_2_2_3_1_2493_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_Minus_2S_2S_1_2495_out1)
          begin :bnn_N_Mux_2_2_3_4_2519
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2519_out1 = bnn_Minus_2S_2S_1_2495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2519_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_Minus_2S_2S_1_2495_out1)
          begin :bnn_N_Mux_2_2_3_1_2520
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2520_out1 = bnn_Minus_2S_2S_1_2495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2520_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1884_out1 or bnn_Minus_2S_2S_1_2468_out1)
          begin :bnn_N_Mux_2_2_3_1_2521
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2521_out1 = bnn_Minus_2S_2S_1_2468_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2521_out1 = bnn_N_Mux_2_2_3_1_1884_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2522
         assign bnn_Minus_2S_2S_1_2522_out1 = -bnn_N_Mux_2_2_3_1_1906_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_6_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4750_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2525_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2525_in2 = {bnn_Mul_16Sx12S_19S_4_4750_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2525_in2 = {{ 5 {fixed_buffer_6_if_1_dout_wire[11]}}, fixed_buffer_6_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2499_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2525_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2525_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2525_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2499_out1[4]}}, bnn_Add_5Sx4S_6S_1_2499_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2525
         assign bnn_Add_17Sx16S_17S_1_2525_out1 = bnn_Add_17Sx16S_17S_1_2525_in2 + {bnn_Add_17Sx16S_17S_1_2525_in1[15], bnn_Add_17Sx16S_17S_1_2525_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2526
         assign bnn_Add_5Sx4S_6S_1_2526_out1 = {bnn_Add_6Ux6U_6U_1_2501_out1[4], bnn_Add_6Ux6U_6U_1_2501_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2500_out1[1]}}, bnn_N_Mux_2_2_3_4_2500_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1941_out1 or bnn_Minus_2S_2S_4_2502_out1)
          begin :bnn_N_Mux_2_2_3_4_2527
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2527_out1 = bnn_Minus_2S_2S_4_2502_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2527_out1 = bnn_N_Mux_2_2_3_1_1941_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2528
         assign bnn_Add_5Sx4S_6S_1_2528_out1 = {bnn_Add_5Sx4S_6S_1_2504_out1[4], bnn_Add_5Sx4S_6S_1_2504_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2503_out1[1]}}, bnn_N_Mux_2_2_3_4_2503_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2529
         assign bnn_Minus_2S_2S_4_2529_out1 = -bnn_N_Mux_2_2_3_1_1952_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1941_out1 or bnn_Minus_2S_2S_4_2502_out1)
          begin :bnn_N_Mux_2_2_3_4_2530
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2530_out1 = bnn_Minus_2S_2S_4_2502_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2530_out1 = bnn_N_Mux_2_2_3_1_1941_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2531
         assign bnn_Add_5Sx4S_6S_1_2531_out1 = {bnn_Add_4Sx2S_5S_1_2507_out1[4], bnn_Add_4Sx2S_5S_1_2507_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2506_out1[1]}}, bnn_N_Mux_2_2_3_4_2506_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1941_out1 or bnn_Minus_2S_2S_4_2502_out1)
          begin :bnn_N_Mux_2_2_3_4_2533
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2533_out1 = bnn_Minus_2S_2S_4_2502_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2533_out1 = bnn_N_Mux_2_2_3_1_1941_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2534
         assign bnn_Add_4Sx2S_5S_1_2534_out1 = {bnn_Add_4Sx2S_4S_1_2510_out1[3], bnn_Add_4Sx2S_4S_1_2510_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2509_out1[1]}}, bnn_N_Mux_2_2_3_4_2509_out1};

         assign bnn_N_Mux_2_2_3_4_2536_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[12], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2511_out1 or bnn_N_Mux_2_2_3_4_2536_in3)
          begin :bnn_N_Mux_2_2_3_4_2536
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2536_out1 = bnn_Minus_2S_2S_4_2511_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2536_out1 = bnn_N_Mux_2_2_3_4_2536_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2537
         assign bnn_Add_4Sx2S_4S_1_2537_out1 = bnn_Add_4Sx2S_4S_1_2513_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2512_out1[1]}}, bnn_N_Mux_2_2_3_4_2512_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2538
         assign bnn_Minus_2S_2S_4_2538_out1 = -bnn_N_Mux_2_4_8_1_1983_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2511_out1 or bnn_N_Mux_2_2_3_4_2536_in3)
          begin :bnn_N_Mux_2_2_3_4_2539
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2539_out1 = bnn_Minus_2S_2S_4_2511_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2539_out1 = bnn_N_Mux_2_2_3_4_2536_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2540
         assign bnn_Add_4Sx2S_4S_1_2540_out1 = bnn_Add_3Sx3S_4S_1_2516_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2515_out1[1]}}, bnn_N_Mux_2_2_3_4_2515_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2511_out1 or bnn_N_Mux_2_2_3_4_2536_in3)
          begin :bnn_N_Mux_2_2_3_4_2542
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2542_out1 = bnn_Minus_2S_2S_4_2511_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2542_out1 = bnn_N_Mux_2_2_3_4_2536_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2543
         assign bnn_Add_3Sx3S_4S_1_2543_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2519_out1[1]}}, bnn_N_Mux_2_2_3_4_2519_out1} + {bnn_Add_2Sx2S_3S_1_2518_out1[2], bnn_Add_2Sx2S_3S_1_2518_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2545
         assign bnn_Add_2Sx2S_3S_1_2545_out1 = {bnn_N_Mux_2_2_3_1_2521_out1[1], bnn_N_Mux_2_2_3_1_2521_out1} + {bnn_N_Mux_2_2_3_1_2520_out1[1], bnn_N_Mux_2_2_3_1_2520_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_Minus_2S_2S_1_2522_out1)
          begin :bnn_N_Mux_2_2_3_4_2546
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2546_out1 = bnn_Minus_2S_2S_1_2522_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2546_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1906_out1 or bnn_Minus_2S_2S_1_2522_out1)
          begin :bnn_N_Mux_2_2_3_1_2547
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2547_out1 = bnn_Minus_2S_2S_1_2522_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2547_out1 = bnn_N_Mux_2_2_3_1_1906_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1895_out1 or bnn_Minus_2S_2S_1_2495_out1)
          begin :bnn_N_Mux_2_2_3_1_2548
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2548_out1 = bnn_Minus_2S_2S_1_2495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2548_out1 = bnn_N_Mux_2_2_3_1_1895_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2549
         assign bnn_Minus_2S_2S_1_2549_out1 = -bnn_N_Mux_2_2_3_1_2158_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2550
         assign bnn_Minus_2S_2S_1_2550_out1 = -bnn_N_Mux_2_2_3_1_1927_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2551
         assign bnn_Minus_2S_2S_1_2551_out1 = -bnn_N_Mux_2_2_3_1_2170_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_7_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4754_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2552_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2552_in2 = {bnn_Mul_16Sx12S_19S_4_4754_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2552_in2 = {{ 5 {fixed_buffer_7_if_1_dout_wire[11]}}, fixed_buffer_7_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2526_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2552_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2552_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2552_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2526_out1[4]}}, bnn_Add_5Sx4S_6S_1_2526_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2552
         assign bnn_Add_17Sx16S_17S_1_2552_out1 = bnn_Add_17Sx16S_17S_1_2552_in2 + {bnn_Add_17Sx16S_17S_1_2552_in1[15], bnn_Add_17Sx16S_17S_1_2552_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2553
         assign bnn_Add_5Sx4S_6S_1_2553_out1 = {bnn_Add_5Sx4S_6S_1_2528_out1[4], bnn_Add_5Sx4S_6S_1_2528_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2527_out1[1]}}, bnn_N_Mux_2_2_3_4_2527_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1952_out1 or bnn_Minus_2S_2S_4_2529_out1)
          begin :bnn_N_Mux_2_2_3_4_2554
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2554_out1 = bnn_Minus_2S_2S_4_2529_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2554_out1 = bnn_N_Mux_2_2_3_1_1952_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2531_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4658_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2555_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2555_in2 = bnn_Mod_5Ux32U_7U_1_4658_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2555_in2 = {bnn_Add_5Sx4S_6S_1_2531_out1[4], bnn_Add_5Sx4S_6S_1_2531_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2530_out1 or bnn_LeftShift_9Ux3U_7U_4_4657_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2555_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2555_in1 = bnn_LeftShift_9Ux3U_7U_4_4657_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2555_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2530_out1[1]}}, bnn_N_Mux_2_2_3_4_2530_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2555
         assign bnn_Add_6Ux6U_6U_1_2555_out1 = bnn_Add_6Ux6U_6U_1_2555_in2 + bnn_Add_6Ux6U_6U_1_2555_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2556
         assign bnn_Minus_2S_2S_4_2556_out1 = -bnn_N_Mux_2_2_3_1_1963_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1952_out1 or bnn_Minus_2S_2S_4_2529_out1)
          begin :bnn_N_Mux_2_2_3_4_2557
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2557_out1 = bnn_Minus_2S_2S_4_2529_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2557_out1 = bnn_N_Mux_2_2_3_1_1952_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2558
         assign bnn_Add_5Sx4S_6S_1_2558_out1 = {bnn_Add_4Sx2S_5S_1_2534_out1[4], bnn_Add_4Sx2S_5S_1_2534_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2533_out1[1]}}, bnn_N_Mux_2_2_3_4_2533_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1952_out1 or bnn_Minus_2S_2S_4_2529_out1)
          begin :bnn_N_Mux_2_2_3_4_2560
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2560_out1 = bnn_Minus_2S_2S_4_2529_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2560_out1 = bnn_N_Mux_2_2_3_1_1952_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2561
         assign bnn_Add_4Sx2S_5S_1_2561_out1 = {bnn_Add_4Sx2S_4S_1_2537_out1[3], bnn_Add_4Sx2S_4S_1_2537_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2536_out1[1]}}, bnn_N_Mux_2_2_3_4_2536_out1};

         assign bnn_N_Mux_2_2_3_4_2563_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[13], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2538_out1 or bnn_N_Mux_2_2_3_4_2563_in3)
          begin :bnn_N_Mux_2_2_3_4_2563
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2563_out1 = bnn_Minus_2S_2S_4_2538_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2563_out1 = bnn_N_Mux_2_2_3_4_2563_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2564
         assign bnn_Add_4Sx2S_4S_1_2564_out1 = bnn_Add_4Sx2S_4S_1_2540_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2539_out1[1]}}, bnn_N_Mux_2_2_3_4_2539_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2565
         assign bnn_Minus_2S_2S_4_2565_out1 = -bnn_N_Mux_2_4_8_1_1994_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2538_out1 or bnn_N_Mux_2_2_3_4_2563_in3)
          begin :bnn_N_Mux_2_2_3_4_2566
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2566_out1 = bnn_Minus_2S_2S_4_2538_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2566_out1 = bnn_N_Mux_2_2_3_4_2563_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2567
         assign bnn_Add_4Sx2S_4S_1_2567_out1 = bnn_Add_3Sx3S_4S_1_2543_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2542_out1[1]}}, bnn_N_Mux_2_2_3_4_2542_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2538_out1 or bnn_N_Mux_2_2_3_4_2563_in3)
          begin :bnn_N_Mux_2_2_3_4_2569
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2569_out1 = bnn_Minus_2S_2S_4_2538_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2569_out1 = bnn_N_Mux_2_2_3_4_2563_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2570
         assign bnn_Add_3Sx3S_4S_1_2570_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2546_out1[1]}}, bnn_N_Mux_2_2_3_4_2546_out1} + {bnn_Add_2Sx2S_3S_1_2545_out1[2], bnn_Add_2Sx2S_3S_1_2545_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2572
         assign bnn_Add_2Sx2S_3S_1_2572_out1 = {bnn_N_Mux_2_2_3_1_2548_out1[1], bnn_N_Mux_2_2_3_1_2548_out1} + {bnn_N_Mux_2_2_3_1_2547_out1[1], bnn_N_Mux_2_2_3_1_2547_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2158_out1 or bnn_Minus_2S_2S_1_2549_out1)
          begin :bnn_N_Mux_2_2_3_4_2573
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2573_out1 = bnn_Minus_2S_2S_1_2549_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2573_out1 = bnn_N_Mux_2_2_3_1_2158_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_Minus_2S_2S_1_2550_out1)
          begin :bnn_N_Mux_2_2_3_4_2574
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2574_out1 = bnn_Minus_2S_2S_1_2550_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2574_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2170_out1 or bnn_Minus_2S_2S_1_2551_out1)
          begin :bnn_N_Mux_2_2_3_4_2575
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2575_out1 = bnn_Minus_2S_2S_1_2551_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2575_out1 = bnn_N_Mux_2_2_3_1_2170_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2576
         assign bnn_Minus_2S_2S_1_2576_out1 = -bnn_N_Mux_2_2_3_1_1938_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_8_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4758_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2579_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2579_in2 = {bnn_Mul_16Sx12S_19S_4_4758_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2579_in2 = {{ 5 {fixed_buffer_8_if_1_dout_wire[11]}}, fixed_buffer_8_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2553_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2579_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2579_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2579_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2553_out1[4]}}, bnn_Add_5Sx4S_6S_1_2553_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2579
         assign bnn_Add_17Sx16S_17S_1_2579_out1 = bnn_Add_17Sx16S_17S_1_2579_in2 + {bnn_Add_17Sx16S_17S_1_2579_in1[15], bnn_Add_17Sx16S_17S_1_2579_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2580
         assign bnn_Add_5Sx4S_6S_1_2580_out1 = {bnn_Add_6Ux6U_6U_1_2555_out1[4], bnn_Add_6Ux6U_6U_1_2555_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2554_out1[1]}}, bnn_N_Mux_2_2_3_4_2554_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1963_out1 or bnn_Minus_2S_2S_4_2556_out1)
          begin :bnn_N_Mux_2_2_3_4_2581
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2581_out1 = bnn_Minus_2S_2S_4_2556_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2581_out1 = bnn_N_Mux_2_2_3_1_1963_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2558_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4667_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2582_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2582_in2 = bnn_Mod_5Ux32U_7U_1_4667_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2582_in2 = {bnn_Add_5Sx4S_6S_1_2558_out1[4], bnn_Add_5Sx4S_6S_1_2558_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2557_out1 or bnn_LeftShift_9Ux3U_7U_4_4666_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2582_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2582_in1 = bnn_LeftShift_9Ux3U_7U_4_4666_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2582_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2557_out1[1]}}, bnn_N_Mux_2_2_3_4_2557_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2582
         assign bnn_Add_6Ux6U_6U_1_2582_out1 = bnn_Add_6Ux6U_6U_1_2582_in2 + bnn_Add_6Ux6U_6U_1_2582_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2583
         assign bnn_Minus_2S_2S_4_2583_out1 = -bnn_N_Mux_2_2_3_1_1974_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1963_out1 or bnn_Minus_2S_2S_4_2556_out1)
          begin :bnn_N_Mux_2_2_3_4_2584
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2584_out1 = bnn_Minus_2S_2S_4_2556_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2584_out1 = bnn_N_Mux_2_2_3_1_1963_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2585
         assign bnn_Add_5Sx4S_6S_1_2585_out1 = {bnn_Add_4Sx2S_5S_1_2561_out1[4], bnn_Add_4Sx2S_5S_1_2561_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2560_out1[1]}}, bnn_N_Mux_2_2_3_4_2560_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1963_out1 or bnn_Minus_2S_2S_4_2556_out1)
          begin :bnn_N_Mux_2_2_3_4_2587
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2587_out1 = bnn_Minus_2S_2S_4_2556_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2587_out1 = bnn_N_Mux_2_2_3_1_1963_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2588
         assign bnn_Add_4Sx2S_5S_1_2588_out1 = {bnn_Add_4Sx2S_4S_1_2564_out1[3], bnn_Add_4Sx2S_4S_1_2564_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2563_out1[1]}}, bnn_N_Mux_2_2_3_4_2563_out1};

         assign bnn_N_Mux_2_2_3_4_2590_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[14], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2565_out1 or bnn_N_Mux_2_2_3_4_2590_in3)
          begin :bnn_N_Mux_2_2_3_4_2590
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2590_out1 = bnn_Minus_2S_2S_4_2565_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2590_out1 = bnn_N_Mux_2_2_3_4_2590_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2591
         assign bnn_Add_4Sx2S_4S_1_2591_out1 = bnn_Add_4Sx2S_4S_1_2567_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2566_out1[1]}}, bnn_N_Mux_2_2_3_4_2566_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2592
         assign bnn_Minus_2S_2S_4_2592_out1 = -bnn_N_Mux_2_4_8_1_2005_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2565_out1 or bnn_N_Mux_2_2_3_4_2590_in3)
          begin :bnn_N_Mux_2_2_3_4_2593
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2593_out1 = bnn_Minus_2S_2S_4_2565_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2593_out1 = bnn_N_Mux_2_2_3_4_2590_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2594
         assign bnn_Add_4Sx2S_4S_1_2594_out1 = bnn_Add_3Sx3S_4S_1_2570_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2569_out1[1]}}, bnn_N_Mux_2_2_3_4_2569_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2565_out1 or bnn_N_Mux_2_2_3_4_2590_in3)
          begin :bnn_N_Mux_2_2_3_4_2596
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2596_out1 = bnn_Minus_2S_2S_4_2565_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2596_out1 = bnn_N_Mux_2_2_3_4_2590_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2597
         assign bnn_Add_3Sx3S_4S_1_2597_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2573_out1[1]}}, bnn_N_Mux_2_2_3_4_2573_out1} + {bnn_Add_2Sx2S_3S_1_2572_out1[2], bnn_Add_2Sx2S_3S_1_2572_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2598
         assign bnn_Minus_2S_2S_4_2598_out1 = -bnn_N_Mux_3_2_6_1_1688_out1_slice;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2599
         assign bnn_Add_2Sx2S_3S_1_2599_out1 = {bnn_N_Mux_2_2_3_4_2575_out1[1], bnn_N_Mux_2_2_3_4_2575_out1} + {bnn_N_Mux_2_2_3_4_2574_out1[1], bnn_N_Mux_2_2_3_4_2574_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_Minus_2S_2S_1_2576_out1)
          begin :bnn_N_Mux_2_2_3_4_2600
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2600_out1 = bnn_Minus_2S_2S_1_2576_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2600_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_Minus_2S_2S_1_2576_out1)
          begin :bnn_N_Mux_2_2_3_1_2601
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_2601_out1 = bnn_Minus_2S_2S_1_2576_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2601_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1927_out1 or bnn_Minus_2S_2S_1_2550_out1)
          begin :bnn_N_Mux_2_2_3_1_2602
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_2602_out1 = bnn_Minus_2S_2S_1_2550_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_2602_out1 = bnn_N_Mux_2_2_3_1_1927_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2603
         assign bnn_Minus_2S_2S_4_2603_out1 = -bnn_N_Mux_2_2_3_1_1949_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_9_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4762_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2606_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2606_in2 = {bnn_Mul_16Sx12S_19S_4_4762_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2606_in2 = {{ 5 {fixed_buffer_9_if_1_dout_wire[11]}}, fixed_buffer_9_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2580_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2606_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2606_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2606_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2580_out1[4]}}, bnn_Add_5Sx4S_6S_1_2580_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2606
         assign bnn_Add_17Sx16S_17S_1_2606_out1 = bnn_Add_17Sx16S_17S_1_2606_in2 + {bnn_Add_17Sx16S_17S_1_2606_in1[15], bnn_Add_17Sx16S_17S_1_2606_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2607
         assign bnn_Add_5Sx4S_6S_1_2607_out1 = {bnn_Add_6Ux6U_6U_1_2582_out1[4], bnn_Add_6Ux6U_6U_1_2582_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2581_out1[1]}}, bnn_N_Mux_2_2_3_4_2581_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1974_out1 or bnn_Minus_2S_2S_4_2583_out1)
          begin :bnn_N_Mux_2_2_3_4_2608
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2608_out1 = bnn_Minus_2S_2S_4_2583_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2608_out1 = bnn_N_Mux_2_2_3_1_1974_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2585_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4676_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2609_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2609_in2 = bnn_Mod_5Ux32U_7U_1_4676_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2609_in2 = {bnn_Add_5Sx4S_6S_1_2585_out1[4], bnn_Add_5Sx4S_6S_1_2585_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2584_out1 or bnn_LeftShift_9Ux3U_7U_4_4675_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2609_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2609_in1 = bnn_LeftShift_9Ux3U_7U_4_4675_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2609_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2584_out1[1]}}, bnn_N_Mux_2_2_3_4_2584_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2609
         assign bnn_Add_6Ux6U_6U_1_2609_out1 = bnn_Add_6Ux6U_6U_1_2609_in2 + bnn_Add_6Ux6U_6U_1_2609_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2610
         assign bnn_Minus_2S_2S_4_2610_out1 = -bnn_N_Mux_2_2_3_1_1985_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1974_out1 or bnn_Minus_2S_2S_4_2583_out1)
          begin :bnn_N_Mux_2_2_3_4_2611
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2611_out1 = bnn_Minus_2S_2S_4_2583_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2611_out1 = bnn_N_Mux_2_2_3_1_1974_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2612
         assign bnn_Add_5Sx4S_6S_1_2612_out1 = {bnn_Add_4Sx2S_5S_1_2588_out1[4], bnn_Add_4Sx2S_5S_1_2588_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2587_out1[1]}}, bnn_N_Mux_2_2_3_4_2587_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1974_out1 or bnn_Minus_2S_2S_4_2583_out1)
          begin :bnn_N_Mux_2_2_3_4_2614
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2614_out1 = bnn_Minus_2S_2S_4_2583_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2614_out1 = bnn_N_Mux_2_2_3_1_1974_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2615
         assign bnn_Add_4Sx2S_5S_1_2615_out1 = {bnn_Add_4Sx2S_4S_1_2591_out1[3], bnn_Add_4Sx2S_4S_1_2591_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2590_out1[1]}}, bnn_N_Mux_2_2_3_4_2590_out1};

         assign bnn_N_Mux_2_2_3_4_2617_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[15], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2592_out1 or bnn_N_Mux_2_2_3_4_2617_in3)
          begin :bnn_N_Mux_2_2_3_4_2617
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2617_out1 = bnn_Minus_2S_2S_4_2592_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2617_out1 = bnn_N_Mux_2_2_3_4_2617_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2618
         assign bnn_Add_4Sx2S_4S_1_2618_out1 = bnn_Add_4Sx2S_4S_1_2594_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2593_out1[1]}}, bnn_N_Mux_2_2_3_4_2593_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2619
         assign bnn_Minus_2S_2S_4_2619_out1 = -bnn_N_Mux_3_2_6_1_1687_out1_slice;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2592_out1 or bnn_N_Mux_2_2_3_4_2617_in3)
          begin :bnn_N_Mux_2_2_3_4_2620
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2620_out1 = bnn_Minus_2S_2S_4_2592_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2620_out1 = bnn_N_Mux_2_2_3_4_2617_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2621
         assign bnn_Add_4Sx2S_4S_1_2621_out1 = bnn_Add_3Sx3S_4S_1_2597_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2596_out1[1]}}, bnn_N_Mux_2_2_3_4_2596_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2622
         assign bnn_Minus_2S_2S_4_2622_out1 = -bnn_N_Mux_2_4_8_1_2016_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2598_out1 or bnn_N_Mux_3_2_6_1_1688_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2623
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2623_out1 = bnn_Minus_2S_2S_4_2598_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2623_out1 = bnn_N_Mux_3_2_6_1_1688_out1_slice;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2624
         assign bnn_Add_3Sx3S_4S_1_2624_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2600_out1[1]}}, bnn_N_Mux_2_2_3_4_2600_out1} + {bnn_Add_2Sx2S_3S_1_2599_out1[2], bnn_Add_2Sx2S_3S_1_2599_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2626
         assign bnn_Add_2Sx2S_3S_1_2626_out1 = {bnn_N_Mux_2_2_3_1_2602_out1[1], bnn_N_Mux_2_2_3_1_2602_out1} + {bnn_N_Mux_2_2_3_1_2601_out1[1], bnn_N_Mux_2_2_3_1_2601_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_Minus_2S_2S_4_2603_out1)
          begin :bnn_N_Mux_2_2_3_4_2627
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2627_out1 = bnn_Minus_2S_2S_4_2603_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2627_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_Minus_2S_2S_4_2603_out1)
          begin :bnn_N_Mux_2_2_3_4_2628
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2628_out1 = bnn_Minus_2S_2S_4_2603_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2628_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1938_out1 or bnn_Minus_2S_2S_1_2576_out1)
          begin :bnn_N_Mux_2_2_3_4_2629
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2629_out1 = bnn_Minus_2S_2S_1_2576_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2629_out1 = bnn_N_Mux_2_2_3_1_1938_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2630
         assign bnn_Minus_2S_2S_4_2630_out1 = -bnn_N_Mux_2_2_3_1_1960_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_10_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4766_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2633_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2633_in2 = {bnn_Mul_16Sx12S_19S_4_4766_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2633_in2 = {{ 5 {fixed_buffer_10_if_1_dout_wire[11]}}, fixed_buffer_10_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2607_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2633_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2633_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2633_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2607_out1[4]}}, bnn_Add_5Sx4S_6S_1_2607_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2633
         assign bnn_Add_17Sx16S_17S_1_2633_out1 = bnn_Add_17Sx16S_17S_1_2633_in2 + {bnn_Add_17Sx16S_17S_1_2633_in1[15], bnn_Add_17Sx16S_17S_1_2633_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2634
         assign bnn_Add_5Sx4S_6S_1_2634_out1 = {bnn_Add_6Ux6U_6U_1_2609_out1[4], bnn_Add_6Ux6U_6U_1_2609_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2608_out1[1]}}, bnn_N_Mux_2_2_3_4_2608_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1985_out1 or bnn_Minus_2S_2S_4_2610_out1)
          begin :bnn_N_Mux_2_2_3_4_2635
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2635_out1 = bnn_Minus_2S_2S_4_2610_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2635_out1 = bnn_N_Mux_2_2_3_1_1985_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2612_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4685_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2636_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2636_in2 = bnn_Mod_5Ux32U_7U_1_4685_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2636_in2 = {bnn_Add_5Sx4S_6S_1_2612_out1[4], bnn_Add_5Sx4S_6S_1_2612_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2611_out1 or bnn_LeftShift_9Ux3U_7U_4_4684_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2636_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2636_in1 = bnn_LeftShift_9Ux3U_7U_4_4684_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2636_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2611_out1[1]}}, bnn_N_Mux_2_2_3_4_2611_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2636
         assign bnn_Add_6Ux6U_6U_1_2636_out1 = bnn_Add_6Ux6U_6U_1_2636_in2 + bnn_Add_6Ux6U_6U_1_2636_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2637
         assign bnn_Minus_2S_2S_4_2637_out1 = -bnn_N_Mux_2_2_3_1_1996_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1985_out1 or bnn_Minus_2S_2S_4_2610_out1)
          begin :bnn_N_Mux_2_2_3_4_2638
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2638_out1 = bnn_Minus_2S_2S_4_2610_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2638_out1 = bnn_N_Mux_2_2_3_1_1985_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2639
         assign bnn_Add_5Sx4S_6S_1_2639_out1 = {bnn_Add_4Sx2S_5S_1_2615_out1[4], bnn_Add_4Sx2S_5S_1_2615_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2614_out1[1]}}, bnn_N_Mux_2_2_3_4_2614_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1985_out1 or bnn_Minus_2S_2S_4_2610_out1)
          begin :bnn_N_Mux_2_2_3_4_2641
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2641_out1 = bnn_Minus_2S_2S_4_2610_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2641_out1 = bnn_N_Mux_2_2_3_1_1985_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2642
         assign bnn_Add_4Sx2S_5S_1_2642_out1 = {bnn_Add_4Sx2S_4S_1_2618_out1[3], bnn_Add_4Sx2S_4S_1_2618_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2617_out1[1]}}, bnn_N_Mux_2_2_3_4_2617_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2619_out1 or bnn_N_Mux_3_2_6_1_1687_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2644
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2644_out1 = bnn_Minus_2S_2S_4_2619_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2644_out1 = bnn_N_Mux_3_2_6_1_1687_out1_slice;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2645
         assign bnn_Add_4Sx2S_4S_1_2645_out1 = bnn_Add_4Sx2S_4S_1_2621_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2620_out1[1]}}, bnn_N_Mux_2_2_3_4_2620_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2646
         assign bnn_Minus_2S_2S_4_2646_out1 = -bnn_N_Mux_2_4_8_1_2033_in3;

         assign bnn_N_Mux_2_2_3_4_2647_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[16], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2622_out1 or bnn_N_Mux_2_2_3_4_2647_in3)
          begin :bnn_N_Mux_2_2_3_4_2647
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2647_out1 = bnn_Minus_2S_2S_4_2622_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2647_out1 = bnn_N_Mux_2_2_3_4_2647_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2648
         assign bnn_Add_4Sx3S_4S_1_2648_out1 = bnn_Add_3Sx3S_4S_1_2624_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2623_out1[1]}}, bnn_N_Mux_2_2_3_4_2623_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2622_out1 or bnn_N_Mux_2_2_3_4_2647_in3)
          begin :bnn_N_Mux_2_2_3_4_2650
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2650_out1 = bnn_Minus_2S_2S_4_2622_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2650_out1 = bnn_N_Mux_2_2_3_4_2647_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2651
         assign bnn_Add_3Sx3S_4S_1_2651_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2627_out1[1]}}, bnn_N_Mux_2_2_3_4_2627_out1} + {bnn_Add_2Sx2S_3S_1_2626_out1[2], bnn_Add_2Sx2S_3S_1_2626_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2653
         assign bnn_Add_2Sx2S_3S_1_2653_out1 = {bnn_N_Mux_2_2_3_4_2629_out1[1], bnn_N_Mux_2_2_3_4_2629_out1} + {bnn_N_Mux_2_2_3_4_2628_out1[1], bnn_N_Mux_2_2_3_4_2628_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_Minus_2S_2S_4_2630_out1)
          begin :bnn_N_Mux_2_2_3_4_2654
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2654_out1 = bnn_Minus_2S_2S_4_2630_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2654_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_Minus_2S_2S_4_2630_out1)
          begin :bnn_N_Mux_2_2_3_4_2655
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2655_out1 = bnn_Minus_2S_2S_4_2630_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2655_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1949_out1 or bnn_Minus_2S_2S_4_2603_out1)
          begin :bnn_N_Mux_2_2_3_4_2656
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2656_out1 = bnn_Minus_2S_2S_4_2603_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2656_out1 = bnn_N_Mux_2_2_3_1_1949_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2657
         assign bnn_Minus_2S_2S_4_2657_out1 = -bnn_N_Mux_2_2_3_1_1971_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_11_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4770_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2660_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2660_in2 = {bnn_Mul_16Sx12S_19S_4_4770_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2660_in2 = {{ 5 {fixed_buffer_11_if_1_dout_wire[11]}}, fixed_buffer_11_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2634_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2660_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2660_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2660_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2634_out1[4]}}, bnn_Add_5Sx4S_6S_1_2634_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2660
         assign bnn_Add_17Sx16S_17S_1_2660_out1 = bnn_Add_17Sx16S_17S_1_2660_in2 + {bnn_Add_17Sx16S_17S_1_2660_in1[15], bnn_Add_17Sx16S_17S_1_2660_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2661
         assign bnn_Add_5Sx4S_6S_1_2661_out1 = {bnn_Add_6Ux6U_6U_1_2636_out1[4], bnn_Add_6Ux6U_6U_1_2636_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2635_out1[1]}}, bnn_N_Mux_2_2_3_4_2635_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1996_out1 or bnn_Minus_2S_2S_4_2637_out1)
          begin :bnn_N_Mux_2_2_3_4_2662
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2662_out1 = bnn_Minus_2S_2S_4_2637_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2662_out1 = bnn_N_Mux_2_2_3_1_1996_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2639_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4694_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2663_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2663_in2 = bnn_Mod_5Ux32U_7U_1_4694_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2663_in2 = {bnn_Add_5Sx4S_6S_1_2639_out1[4], bnn_Add_5Sx4S_6S_1_2639_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2638_out1 or bnn_LeftShift_9Ux3U_7U_4_4693_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2663_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2663_in1 = bnn_LeftShift_9Ux3U_7U_4_4693_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2663_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2638_out1[1]}}, bnn_N_Mux_2_2_3_4_2638_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2663
         assign bnn_Add_6Ux6U_6U_1_2663_out1 = bnn_Add_6Ux6U_6U_1_2663_in2 + bnn_Add_6Ux6U_6U_1_2663_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2664
         assign bnn_Minus_2S_2S_4_2664_out1 = -bnn_N_Mux_2_2_3_1_2007_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1996_out1 or bnn_Minus_2S_2S_4_2637_out1)
          begin :bnn_N_Mux_2_2_3_4_2665
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2665_out1 = bnn_Minus_2S_2S_4_2637_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2665_out1 = bnn_N_Mux_2_2_3_1_1996_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2666
         assign bnn_Add_5Sx4S_6S_1_2666_out1 = {bnn_Add_4Sx2S_5S_1_2642_out1[4], bnn_Add_4Sx2S_5S_1_2642_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2641_out1[1]}}, bnn_N_Mux_2_2_3_4_2641_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1996_out1 or bnn_Minus_2S_2S_4_2637_out1)
          begin :bnn_N_Mux_2_2_3_4_2668
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2668_out1 = bnn_Minus_2S_2S_4_2637_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2668_out1 = bnn_N_Mux_2_2_3_1_1996_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2669
         assign bnn_Add_4Sx2S_5S_1_2669_out1 = {bnn_Add_4Sx2S_4S_1_2645_out1[3], bnn_Add_4Sx2S_4S_1_2645_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2644_out1[1]}}, bnn_N_Mux_2_2_3_4_2644_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2670
         assign bnn_Minus_2S_2S_4_2670_out1 = -bnn_N_Mux_2_2_3_1_2205_out1;

         assign bnn_N_Mux_2_2_3_4_2671_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[17], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2646_out1 or bnn_N_Mux_2_2_3_4_2671_in3)
          begin :bnn_N_Mux_2_2_3_4_2671
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2671_out1 = bnn_Minus_2S_2S_4_2646_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2671_out1 = bnn_N_Mux_2_2_3_4_2671_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2672
         assign bnn_Add_4Sx3S_4S_1_2672_out1 = bnn_Add_4Sx3S_4S_1_2648_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2647_out1[1]}}, bnn_N_Mux_2_2_3_4_2647_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2673
         assign bnn_Minus_2S_2S_4_2673_out1 = -bnn_N_Mux_2_4_8_1_2050_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2646_out1 or bnn_N_Mux_2_2_3_4_2671_in3)
          begin :bnn_N_Mux_2_2_3_4_2674
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2674_out1 = bnn_Minus_2S_2S_4_2646_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2674_out1 = bnn_N_Mux_2_2_3_4_2671_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2675
         assign bnn_Add_4Sx2S_4S_1_2675_out1 = bnn_Add_3Sx3S_4S_1_2651_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2650_out1[1]}}, bnn_N_Mux_2_2_3_4_2650_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2646_out1 or bnn_N_Mux_2_2_3_4_2671_in3)
          begin :bnn_N_Mux_2_2_3_4_2677
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2677_out1 = bnn_Minus_2S_2S_4_2646_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2677_out1 = bnn_N_Mux_2_2_3_4_2671_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2678
         assign bnn_Add_3Sx3S_4S_1_2678_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2654_out1[1]}}, bnn_N_Mux_2_2_3_4_2654_out1} + {bnn_Add_2Sx2S_3S_1_2653_out1[2], bnn_Add_2Sx2S_3S_1_2653_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2680
         assign bnn_Add_2Sx2S_3S_1_2680_out1 = {bnn_N_Mux_2_2_3_4_2656_out1[1], bnn_N_Mux_2_2_3_4_2656_out1} + {bnn_N_Mux_2_2_3_4_2655_out1[1], bnn_N_Mux_2_2_3_4_2655_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_Minus_2S_2S_4_2657_out1)
          begin :bnn_N_Mux_2_2_3_4_2681
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2681_out1 = bnn_Minus_2S_2S_4_2657_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2681_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_Minus_2S_2S_4_2657_out1)
          begin :bnn_N_Mux_2_2_3_4_2682
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2682_out1 = bnn_Minus_2S_2S_4_2657_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2682_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1960_out1 or bnn_Minus_2S_2S_4_2630_out1)
          begin :bnn_N_Mux_2_2_3_4_2683
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2683_out1 = bnn_Minus_2S_2S_4_2630_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2683_out1 = bnn_N_Mux_2_2_3_1_1960_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2684
         assign bnn_Minus_2S_2S_4_2684_out1 = -bnn_N_Mux_2_2_3_1_1982_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_12_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4774_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2687_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2687_in2 = {bnn_Mul_16Sx12S_19S_4_4774_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2687_in2 = {{ 5 {fixed_buffer_12_if_1_dout_wire[11]}}, fixed_buffer_12_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2661_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2687_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2687_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2687_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2661_out1[4]}}, bnn_Add_5Sx4S_6S_1_2661_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2687
         assign bnn_Add_17Sx16S_17S_1_2687_out1 = bnn_Add_17Sx16S_17S_1_2687_in2 + {bnn_Add_17Sx16S_17S_1_2687_in1[15], bnn_Add_17Sx16S_17S_1_2687_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2688
         assign bnn_Add_5Sx4S_6S_1_2688_out1 = {bnn_Add_6Ux6U_6U_1_2663_out1[4], bnn_Add_6Ux6U_6U_1_2663_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2662_out1[1]}}, bnn_N_Mux_2_2_3_4_2662_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2007_out1 or bnn_Minus_2S_2S_4_2664_out1)
          begin :bnn_N_Mux_2_2_3_4_2689
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2689_out1 = bnn_Minus_2S_2S_4_2664_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2689_out1 = bnn_N_Mux_2_2_3_1_2007_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2666_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4703_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2690_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2690_in2 = bnn_Mod_5Ux32U_7U_1_4703_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2690_in2 = {bnn_Add_5Sx4S_6S_1_2666_out1[4], bnn_Add_5Sx4S_6S_1_2666_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2665_out1 or bnn_LeftShift_9Ux3U_7U_4_4702_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2690_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2690_in1 = bnn_LeftShift_9Ux3U_7U_4_4702_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2690_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2665_out1[1]}}, bnn_N_Mux_2_2_3_4_2665_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2690
         assign bnn_Add_6Ux6U_6U_1_2690_out1 = bnn_Add_6Ux6U_6U_1_2690_in2 + bnn_Add_6Ux6U_6U_1_2690_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2691
         assign bnn_Minus_2S_2S_4_2691_out1 = -bnn_N_Mux_2_2_3_1_2187_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2007_out1 or bnn_Minus_2S_2S_4_2664_out1)
          begin :bnn_N_Mux_2_2_3_4_2692
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2692_out1 = bnn_Minus_2S_2S_4_2664_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2692_out1 = bnn_N_Mux_2_2_3_1_2007_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2693
         assign bnn_Add_5Sx4S_6S_1_2693_out1 = {bnn_Add_4Sx2S_5S_1_2669_out1[4], bnn_Add_4Sx2S_5S_1_2669_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2668_out1[1]}}, bnn_N_Mux_2_2_3_4_2668_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2694
         assign bnn_Minus_2S_2S_4_2694_out1 = -bnn_N_Mux_2_2_3_1_2018_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2205_out1 or bnn_Minus_2S_2S_4_2670_out1)
          begin :bnn_N_Mux_2_2_3_4_2695
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2695_out1 = bnn_Minus_2S_2S_4_2670_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2695_out1 = bnn_N_Mux_2_2_3_1_2205_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2696
         assign bnn_Add_4Sx2S_5S_1_2696_out1 = {bnn_Add_4Sx3S_4S_1_2672_out1[3], bnn_Add_4Sx3S_4S_1_2672_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2671_out1[1]}}, bnn_N_Mux_2_2_3_4_2671_out1};

         assign bnn_N_Mux_2_2_3_4_2698_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[18], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2673_out1 or bnn_N_Mux_2_2_3_4_2698_in3)
          begin :bnn_N_Mux_2_2_3_4_2698
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2698_out1 = bnn_Minus_2S_2S_4_2673_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2698_out1 = bnn_N_Mux_2_2_3_4_2698_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_2699
         assign bnn_Add_4Sx2S_4S_1_2699_out1 = bnn_Add_4Sx2S_4S_1_2675_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2674_out1[1]}}, bnn_N_Mux_2_2_3_4_2674_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2700
         assign bnn_Minus_2S_2S_4_2700_out1 = -bnn_N_Mux_2_4_8_1_2067_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2673_out1 or bnn_N_Mux_2_2_3_4_2698_in3)
          begin :bnn_N_Mux_2_2_3_4_2701
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2701_out1 = bnn_Minus_2S_2S_4_2673_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2701_out1 = bnn_N_Mux_2_2_3_4_2698_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2702
         assign bnn_Add_4Sx3S_4S_1_2702_out1 = bnn_Add_3Sx3S_4S_1_2678_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2677_out1[1]}}, bnn_N_Mux_2_2_3_4_2677_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2673_out1 or bnn_N_Mux_2_2_3_4_2698_in3)
          begin :bnn_N_Mux_2_2_3_4_2704
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2704_out1 = bnn_Minus_2S_2S_4_2673_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2704_out1 = bnn_N_Mux_2_2_3_4_2698_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2705
         assign bnn_Add_3Sx3S_4S_1_2705_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2681_out1[1]}}, bnn_N_Mux_2_2_3_4_2681_out1} + {bnn_Add_2Sx2S_3S_1_2680_out1[2], bnn_Add_2Sx2S_3S_1_2680_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2707
         assign bnn_Add_2Sx2S_3S_1_2707_out1 = {bnn_N_Mux_2_2_3_4_2683_out1[1], bnn_N_Mux_2_2_3_4_2683_out1} + {bnn_N_Mux_2_2_3_4_2682_out1[1], bnn_N_Mux_2_2_3_4_2682_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_Minus_2S_2S_4_2684_out1)
          begin :bnn_N_Mux_2_2_3_4_2708
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2708_out1 = bnn_Minus_2S_2S_4_2684_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2708_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_Minus_2S_2S_4_2684_out1)
          begin :bnn_N_Mux_2_2_3_4_2709
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2709_out1 = bnn_Minus_2S_2S_4_2684_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2709_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1971_out1 or bnn_Minus_2S_2S_4_2657_out1)
          begin :bnn_N_Mux_2_2_3_4_2710
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2710_out1 = bnn_Minus_2S_2S_4_2657_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2710_out1 = bnn_N_Mux_2_2_3_1_1971_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2711
         assign bnn_Minus_2S_2S_4_2711_out1 = -bnn_N_Mux_2_2_3_1_1993_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_13_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4778_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2714_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2714_in2 = {bnn_Mul_16Sx12S_19S_4_4778_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2714_in2 = {{ 5 {fixed_buffer_13_if_1_dout_wire[11]}}, fixed_buffer_13_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2688_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2714_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2714_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2714_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2688_out1[4]}}, bnn_Add_5Sx4S_6S_1_2688_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2714
         assign bnn_Add_17Sx16S_17S_1_2714_out1 = bnn_Add_17Sx16S_17S_1_2714_in2 + {bnn_Add_17Sx16S_17S_1_2714_in1[15], bnn_Add_17Sx16S_17S_1_2714_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2715
         assign bnn_Add_5Sx4S_6S_1_2715_out1 = {bnn_Add_6Ux6U_6U_1_2690_out1[4], bnn_Add_6Ux6U_6U_1_2690_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2689_out1[1]}}, bnn_N_Mux_2_2_3_4_2689_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2187_out1 or bnn_Minus_2S_2S_4_2691_out1)
          begin :bnn_N_Mux_2_2_3_4_2716
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2716_out1 = bnn_Minus_2S_2S_4_2691_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2716_out1 = bnn_N_Mux_2_2_3_1_2187_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2693_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4712_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2717_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2717_in2 = bnn_Mod_5Ux32U_7U_1_4712_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2717_in2 = {bnn_Add_5Sx4S_6S_1_2693_out1[4], bnn_Add_5Sx4S_6S_1_2693_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2692_out1 or bnn_LeftShift_9Ux3U_7U_4_4711_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2717_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2717_in1 = bnn_LeftShift_9Ux3U_7U_4_4711_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2717_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2692_out1[1]}}, bnn_N_Mux_2_2_3_4_2692_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2717
         assign bnn_Add_6Ux6U_6U_1_2717_out1 = bnn_Add_6Ux6U_6U_1_2717_in2 + bnn_Add_6Ux6U_6U_1_2717_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2718
         assign bnn_Minus_2S_2S_4_2718_out1 = -bnn_N_Mux_2_2_3_1_2035_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2018_out1 or bnn_Minus_2S_2S_4_2694_out1)
          begin :bnn_N_Mux_2_2_3_4_2719
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2719_out1 = bnn_Minus_2S_2S_4_2694_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2719_out1 = bnn_N_Mux_2_2_3_1_2018_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2720
         assign bnn_Add_5Sx4S_6S_1_2720_out1 = {bnn_Add_4Sx2S_5S_1_2696_out1[4], bnn_Add_4Sx2S_5S_1_2696_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2695_out1[1]}}, bnn_N_Mux_2_2_3_4_2695_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2018_out1 or bnn_Minus_2S_2S_4_2694_out1)
          begin :bnn_N_Mux_2_2_3_4_2722
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2722_out1 = bnn_Minus_2S_2S_4_2694_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2722_out1 = bnn_N_Mux_2_2_3_1_2018_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2723
         assign bnn_Add_4Sx2S_5S_1_2723_out1 = {bnn_Add_4Sx2S_4S_1_2699_out1[3], bnn_Add_4Sx2S_4S_1_2699_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2698_out1[1]}}, bnn_N_Mux_2_2_3_4_2698_out1};

         assign bnn_N_Mux_2_2_3_4_2725_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[19], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2700_out1 or bnn_N_Mux_2_2_3_4_2725_in3)
          begin :bnn_N_Mux_2_2_3_4_2725
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2725_out1 = bnn_Minus_2S_2S_4_2700_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2725_out1 = bnn_N_Mux_2_2_3_4_2725_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2726
         assign bnn_Add_4Sx3S_4S_1_2726_out1 = bnn_Add_4Sx3S_4S_1_2702_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2701_out1[1]}}, bnn_N_Mux_2_2_3_4_2701_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2727
         assign bnn_Minus_2S_2S_4_2727_out1 = -bnn_N_Mux_2_4_8_1_2084_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2700_out1 or bnn_N_Mux_2_2_3_4_2725_in3)
          begin :bnn_N_Mux_2_2_3_4_2728
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2728_out1 = bnn_Minus_2S_2S_4_2700_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2728_out1 = bnn_N_Mux_2_2_3_4_2725_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2729
         assign bnn_Add_4Sx3S_4S_1_2729_out1 = bnn_Add_3Sx3S_4S_1_2705_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2704_out1[1]}}, bnn_N_Mux_2_2_3_4_2704_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2700_out1 or bnn_N_Mux_2_2_3_4_2725_in3)
          begin :bnn_N_Mux_2_2_3_4_2731
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2731_out1 = bnn_Minus_2S_2S_4_2700_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2731_out1 = bnn_N_Mux_2_2_3_4_2725_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2732
         assign bnn_Add_3Sx3S_4S_1_2732_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2708_out1[1]}}, bnn_N_Mux_2_2_3_4_2708_out1} + {bnn_Add_2Sx2S_3S_1_2707_out1[2], bnn_Add_2Sx2S_3S_1_2707_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2734
         assign bnn_Add_2Sx2S_3S_1_2734_out1 = {bnn_N_Mux_2_2_3_4_2710_out1[1], bnn_N_Mux_2_2_3_4_2710_out1} + {bnn_N_Mux_2_2_3_4_2709_out1[1], bnn_N_Mux_2_2_3_4_2709_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_Minus_2S_2S_4_2711_out1)
          begin :bnn_N_Mux_2_2_3_4_2735
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2735_out1 = bnn_Minus_2S_2S_4_2711_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2735_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_Minus_2S_2S_4_2711_out1)
          begin :bnn_N_Mux_2_2_3_4_2736
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2736_out1 = bnn_Minus_2S_2S_4_2711_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2736_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1982_out1 or bnn_Minus_2S_2S_4_2684_out1)
          begin :bnn_N_Mux_2_2_3_4_2737
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2737_out1 = bnn_Minus_2S_2S_4_2684_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2737_out1 = bnn_N_Mux_2_2_3_1_1982_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2738
         assign bnn_Minus_2S_2S_4_2738_out1 = -bnn_N_Mux_2_2_3_1_2004_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_14_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4782_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2741_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2741_in2 = {bnn_Mul_16Sx12S_19S_4_4782_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2741_in2 = {{ 5 {fixed_buffer_14_if_1_dout_wire[11]}}, fixed_buffer_14_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2715_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2741_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2741_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2741_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2715_out1[4]}}, bnn_Add_5Sx4S_6S_1_2715_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2741
         assign bnn_Add_17Sx16S_17S_1_2741_out1 = bnn_Add_17Sx16S_17S_1_2741_in2 + {bnn_Add_17Sx16S_17S_1_2741_in1[15], bnn_Add_17Sx16S_17S_1_2741_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2742
         assign bnn_Add_5Sx4S_6S_1_2742_out1 = {bnn_Add_6Ux6U_6U_1_2717_out1[4], bnn_Add_6Ux6U_6U_1_2717_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2716_out1[1]}}, bnn_N_Mux_2_2_3_4_2716_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2035_out1 or bnn_Minus_2S_2S_4_2718_out1)
          begin :bnn_N_Mux_2_2_3_4_2743
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2743_out1 = bnn_Minus_2S_2S_4_2718_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2743_out1 = bnn_N_Mux_2_2_3_1_2035_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2744
         assign bnn_Add_5Sx4S_6S_1_2744_out1 = {bnn_Add_5Sx4S_6S_1_2720_out1[4], bnn_Add_5Sx4S_6S_1_2720_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2719_out1[1]}}, bnn_N_Mux_2_2_3_4_2719_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2745
         assign bnn_Minus_2S_2S_4_2745_out1 = -bnn_N_Mux_2_2_3_1_2052_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2035_out1 or bnn_Minus_2S_2S_4_2718_out1)
          begin :bnn_N_Mux_2_2_3_4_2746
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2746_out1 = bnn_Minus_2S_2S_4_2718_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2746_out1 = bnn_N_Mux_2_2_3_1_2035_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2747
         assign bnn_Add_5Sx4S_6S_1_2747_out1 = {bnn_Add_4Sx2S_5S_1_2723_out1[4], bnn_Add_4Sx2S_5S_1_2723_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2722_out1[1]}}, bnn_N_Mux_2_2_3_4_2722_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2035_out1 or bnn_Minus_2S_2S_4_2718_out1)
          begin :bnn_N_Mux_2_2_3_4_2749
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2749_out1 = bnn_Minus_2S_2S_4_2718_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2749_out1 = bnn_N_Mux_2_2_3_1_2035_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2750
         assign bnn_Add_4Sx2S_5S_1_2750_out1 = {bnn_Add_4Sx3S_4S_1_2726_out1[3], bnn_Add_4Sx3S_4S_1_2726_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2725_out1[1]}}, bnn_N_Mux_2_2_3_4_2725_out1};

         assign bnn_N_Mux_2_2_3_4_2752_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[20], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2727_out1 or bnn_N_Mux_2_2_3_4_2752_in3)
          begin :bnn_N_Mux_2_2_3_4_2752
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2752_out1 = bnn_Minus_2S_2S_4_2727_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2752_out1 = bnn_N_Mux_2_2_3_4_2752_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2753
         assign bnn_Add_4Sx3S_4S_1_2753_out1 = bnn_Add_4Sx3S_4S_1_2729_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2728_out1[1]}}, bnn_N_Mux_2_2_3_4_2728_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2754
         assign bnn_Minus_2S_2S_4_2754_out1 = -bnn_N_Mux_2_4_8_1_2101_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2727_out1 or bnn_N_Mux_2_2_3_4_2752_in3)
          begin :bnn_N_Mux_2_2_3_4_2755
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2755_out1 = bnn_Minus_2S_2S_4_2727_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2755_out1 = bnn_N_Mux_2_2_3_4_2752_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2756
         assign bnn_Add_4Sx3S_4S_1_2756_out1 = bnn_Add_3Sx3S_4S_1_2732_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2731_out1[1]}}, bnn_N_Mux_2_2_3_4_2731_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2727_out1 or bnn_N_Mux_2_2_3_4_2752_in3)
          begin :bnn_N_Mux_2_2_3_4_2758
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2758_out1 = bnn_Minus_2S_2S_4_2727_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2758_out1 = bnn_N_Mux_2_2_3_4_2752_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2759
         assign bnn_Add_3Sx3S_4S_1_2759_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2735_out1[1]}}, bnn_N_Mux_2_2_3_4_2735_out1} + {bnn_Add_2Sx2S_3S_1_2734_out1[2], bnn_Add_2Sx2S_3S_1_2734_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2761
         assign bnn_Add_2Sx2S_3S_1_2761_out1 = {bnn_N_Mux_2_2_3_4_2737_out1[1], bnn_N_Mux_2_2_3_4_2737_out1} + {bnn_N_Mux_2_2_3_4_2736_out1[1], bnn_N_Mux_2_2_3_4_2736_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_Minus_2S_2S_4_2738_out1)
          begin :bnn_N_Mux_2_2_3_4_2762
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2762_out1 = bnn_Minus_2S_2S_4_2738_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2762_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2004_out1 or bnn_Minus_2S_2S_4_2738_out1)
          begin :bnn_N_Mux_2_2_3_4_2763
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2763_out1 = bnn_Minus_2S_2S_4_2738_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2763_out1 = bnn_N_Mux_2_2_3_1_2004_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_1993_out1 or bnn_Minus_2S_2S_4_2711_out1)
          begin :bnn_N_Mux_2_2_3_4_2764
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2764_out1 = bnn_Minus_2S_2S_4_2711_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2764_out1 = bnn_N_Mux_2_2_3_1_1993_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2765
         assign bnn_Minus_2S_2S_4_2765_out1 = -bnn_N_Mux_2_2_3_1_2184_out1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2766
         assign bnn_Minus_2S_2S_4_2766_out1 = -bnn_N_Mux_2_2_3_1_2015_out1;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2767
         assign bnn_Minus_2S_2S_1_2767_out1 = -bnn_N_Mux_2_2_3_1_2202_out1;

         assign bnn_N_Mux_3_2_6_4_2768_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[23], bnn_N_Mux_64_2_2_1_1636_out1[23]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_2768_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_2768
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_2768_out1_slice = bnn_N_Mux_3_2_6_4_2768_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_2768_out1_slice = 2'd0;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_15_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4786_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2769_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2769_in2 = {bnn_Mul_16Sx12S_19S_4_4786_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2769_in2 = {{ 5 {fixed_buffer_15_if_1_dout_wire[11]}}, fixed_buffer_15_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2742_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2769_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2769_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2769_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2742_out1[4]}}, bnn_Add_5Sx4S_6S_1_2742_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2769
         assign bnn_Add_17Sx16S_17S_1_2769_out1 = bnn_Add_17Sx16S_17S_1_2769_in2 + {bnn_Add_17Sx16S_17S_1_2769_in1[15], bnn_Add_17Sx16S_17S_1_2769_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2770
         assign bnn_Add_5Sx4S_6S_1_2770_out1 = {bnn_Add_5Sx4S_6S_1_2744_out1[4], bnn_Add_5Sx4S_6S_1_2744_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2743_out1[1]}}, bnn_N_Mux_2_2_3_4_2743_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2052_out1 or bnn_Minus_2S_2S_4_2745_out1)
          begin :bnn_N_Mux_2_2_3_4_2771
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2771_out1 = bnn_Minus_2S_2S_4_2745_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2771_out1 = bnn_N_Mux_2_2_3_1_2052_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_2747_out1[4:0] or bnn_Mod_5Ux32U_7U_1_4721_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2772_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2772_in2 = bnn_Mod_5Ux32U_7U_1_4721_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2772_in2 = {bnn_Add_5Sx4S_6S_1_2747_out1[4], bnn_Add_5Sx4S_6S_1_2747_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(bnn_N_Mux_2_2_3_4_2746_out1 or bnn_LeftShift_9Ux3U_7U_4_4720_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_2772_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_2772_in1 = bnn_LeftShift_9Ux3U_7U_4_4720_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_2772_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_2746_out1[1]}}, bnn_N_Mux_2_2_3_4_2746_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_2772
         assign bnn_Add_6Ux6U_6U_1_2772_out1 = bnn_Add_6Ux6U_6U_1_2772_in2 + bnn_Add_6Ux6U_6U_1_2772_in1;

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2773
         assign bnn_Minus_2S_2S_4_2773_out1 = -bnn_N_Mux_2_2_3_1_2069_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2052_out1 or bnn_Minus_2S_2S_4_2745_out1)
          begin :bnn_N_Mux_2_2_3_4_2774
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2774_out1 = bnn_Minus_2S_2S_4_2745_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2774_out1 = bnn_N_Mux_2_2_3_1_2052_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2775
         assign bnn_Add_5Sx4S_6S_1_2775_out1 = {bnn_Add_4Sx2S_5S_1_2750_out1[4], bnn_Add_4Sx2S_5S_1_2750_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2749_out1[1]}}, bnn_N_Mux_2_2_3_4_2749_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2052_out1 or bnn_Minus_2S_2S_4_2745_out1)
          begin :bnn_N_Mux_2_2_3_4_2777
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2777_out1 = bnn_Minus_2S_2S_4_2745_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2777_out1 = bnn_N_Mux_2_2_3_1_2052_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2778
         assign bnn_Add_4Sx2S_5S_1_2778_out1 = {bnn_Add_4Sx3S_4S_1_2753_out1[3], bnn_Add_4Sx3S_4S_1_2753_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2752_out1[1]}}, bnn_N_Mux_2_2_3_4_2752_out1};

         assign bnn_N_Mux_2_2_3_4_2780_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[21], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2754_out1 or bnn_N_Mux_2_2_3_4_2780_in3)
          begin :bnn_N_Mux_2_2_3_4_2780
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2780_out1 = bnn_Minus_2S_2S_4_2754_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2780_out1 = bnn_N_Mux_2_2_3_4_2780_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2781
         assign bnn_Add_4Sx3S_4S_1_2781_out1 = bnn_Add_4Sx3S_4S_1_2756_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2755_out1[1]}}, bnn_N_Mux_2_2_3_4_2755_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2782
         assign bnn_Minus_2S_2S_4_2782_out1 = -bnn_N_Mux_2_4_8_1_2118_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2754_out1 or bnn_N_Mux_2_2_3_4_2780_in3)
          begin :bnn_N_Mux_2_2_3_4_2783
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2783_out1 = bnn_Minus_2S_2S_4_2754_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2783_out1 = bnn_N_Mux_2_2_3_4_2780_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2784
         assign bnn_Add_4Sx3S_4S_1_2784_out1 = bnn_Add_3Sx3S_4S_1_2759_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2758_out1[1]}}, bnn_N_Mux_2_2_3_4_2758_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2754_out1 or bnn_N_Mux_2_2_3_4_2780_in3)
          begin :bnn_N_Mux_2_2_3_4_2786
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2786_out1 = bnn_Minus_2S_2S_4_2754_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2786_out1 = bnn_N_Mux_2_2_3_4_2780_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2787
         assign bnn_Add_3Sx3S_4S_1_2787_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2762_out1[1]}}, bnn_N_Mux_2_2_3_4_2762_out1} + {bnn_Add_2Sx2S_3S_1_2761_out1[2], bnn_Add_2Sx2S_3S_1_2761_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2789
         assign bnn_Add_2Sx2S_3S_1_2789_out1 = {bnn_N_Mux_2_2_3_4_2764_out1[1], bnn_N_Mux_2_2_3_4_2764_out1} + {bnn_N_Mux_2_2_3_4_2763_out1[1], bnn_N_Mux_2_2_3_4_2763_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2184_out1 or bnn_Minus_2S_2S_4_2765_out1)
          begin :bnn_N_Mux_2_2_3_4_2790
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2790_out1 = bnn_Minus_2S_2S_4_2765_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2790_out1 = bnn_N_Mux_2_2_3_1_2184_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_Minus_2S_2S_4_2766_out1)
          begin :bnn_N_Mux_2_2_3_4_2791
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2791_out1 = bnn_Minus_2S_2S_4_2766_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2791_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2202_out1 or bnn_Minus_2S_2S_1_2767_out1)
          begin :bnn_N_Mux_2_2_3_4_2792
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2792_out1 = bnn_Minus_2S_2S_1_2767_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2792_out1 = bnn_N_Mux_2_2_3_1_2202_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2793
         assign bnn_Minus_2S_2S_4_2793_out1 = -bnn_N_Mux_2_2_3_1_2032_out1;

         assign bnn_N_Mux_3_2_6_4_2796_in2 = {{bnn_N_Mux_64_2_2_1_1636_out1[24], bnn_N_Mux_64_2_2_1_1636_out1[24]}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_2796_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_2796
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_2796_out1_slice = bnn_N_Mux_3_2_6_4_2796_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_2796_out1_slice = 2'd0;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_16_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4790_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2797_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2797_in2 = {bnn_Mul_16Sx12S_19S_4_4790_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2797_in2 = {{ 5 {fixed_buffer_16_if_1_dout_wire[11]}}, fixed_buffer_16_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2770_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2797_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2797_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2797_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2770_out1[4]}}, bnn_Add_5Sx4S_6S_1_2770_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2797
         assign bnn_Add_17Sx16S_17S_1_2797_out1 = bnn_Add_17Sx16S_17S_1_2797_in2 + {bnn_Add_17Sx16S_17S_1_2797_in1[15], bnn_Add_17Sx16S_17S_1_2797_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2798
         assign bnn_Add_5Sx4S_6S_1_2798_out1 = {bnn_Add_6Ux6U_6U_1_2772_out1[4], bnn_Add_6Ux6U_6U_1_2772_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2771_out1[1]}}, bnn_N_Mux_2_2_3_4_2771_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2069_out1 or bnn_Minus_2S_2S_4_2773_out1)
          begin :bnn_N_Mux_2_2_3_4_2799
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2799_out1 = bnn_Minus_2S_2S_4_2773_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2799_out1 = bnn_N_Mux_2_2_3_1_2069_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2800
         assign bnn_Add_5Sx4S_6S_1_2800_out1 = {bnn_Add_5Sx4S_6S_1_2775_out1[4], bnn_Add_5Sx4S_6S_1_2775_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2774_out1[1]}}, bnn_N_Mux_2_2_3_4_2774_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2801
         assign bnn_Minus_2S_2S_4_2801_out1 = -bnn_N_Mux_2_2_3_1_2086_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2069_out1 or bnn_Minus_2S_2S_4_2773_out1)
          begin :bnn_N_Mux_2_2_3_4_2802
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2802_out1 = bnn_Minus_2S_2S_4_2773_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2802_out1 = bnn_N_Mux_2_2_3_1_2069_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2803
         assign bnn_Add_5Sx4S_6S_1_2803_out1 = {bnn_Add_4Sx2S_5S_1_2778_out1[4], bnn_Add_4Sx2S_5S_1_2778_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2777_out1[1]}}, bnn_N_Mux_2_2_3_4_2777_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2069_out1 or bnn_Minus_2S_2S_4_2773_out1)
          begin :bnn_N_Mux_2_2_3_4_2805
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2805_out1 = bnn_Minus_2S_2S_4_2773_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2805_out1 = bnn_N_Mux_2_2_3_1_2069_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2806
         assign bnn_Add_4Sx2S_5S_1_2806_out1 = {bnn_Add_4Sx3S_4S_1_2781_out1[3], bnn_Add_4Sx3S_4S_1_2781_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2780_out1[1]}}, bnn_N_Mux_2_2_3_4_2780_out1};

         assign bnn_N_Mux_2_2_3_4_2808_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[22], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2782_out1 or bnn_N_Mux_2_2_3_4_2808_in3)
          begin :bnn_N_Mux_2_2_3_4_2808
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2808_out1 = bnn_Minus_2S_2S_4_2782_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2808_out1 = bnn_N_Mux_2_2_3_4_2808_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2809
         assign bnn_Add_4Sx3S_4S_1_2809_out1 = bnn_Add_4Sx3S_4S_1_2784_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2783_out1[1]}}, bnn_N_Mux_2_2_3_4_2783_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2810
         assign bnn_Minus_2S_2S_4_2810_out1 = -bnn_N_Mux_2_4_8_1_2135_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2782_out1 or bnn_N_Mux_2_2_3_4_2808_in3)
          begin :bnn_N_Mux_2_2_3_4_2811
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2811_out1 = bnn_Minus_2S_2S_4_2782_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2811_out1 = bnn_N_Mux_2_2_3_4_2808_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2812
         assign bnn_Add_4Sx3S_4S_1_2812_out1 = bnn_Add_3Sx3S_4S_1_2787_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2786_out1[1]}}, bnn_N_Mux_2_2_3_4_2786_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2782_out1 or bnn_N_Mux_2_2_3_4_2808_in3)
          begin :bnn_N_Mux_2_2_3_4_2814
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2814_out1 = bnn_Minus_2S_2S_4_2782_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2814_out1 = bnn_N_Mux_2_2_3_4_2808_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2815
         assign bnn_Add_3Sx3S_4S_1_2815_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2790_out1[1]}}, bnn_N_Mux_2_2_3_4_2790_out1} + {bnn_Add_2Sx2S_3S_1_2789_out1[2], bnn_Add_2Sx2S_3S_1_2789_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2816
         assign bnn_Minus_2S_2S_4_2816_out1 = -bnn_N_Mux_3_2_6_4_2768_out1_slice;

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2817
         assign bnn_Add_2Sx2S_3S_1_2817_out1 = {bnn_N_Mux_2_2_3_4_2792_out1[1], bnn_N_Mux_2_2_3_4_2792_out1} + {bnn_N_Mux_2_2_3_4_2791_out1[1], bnn_N_Mux_2_2_3_4_2791_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_Minus_2S_2S_4_2793_out1)
          begin :bnn_N_Mux_2_2_3_4_2818
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2818_out1 = bnn_Minus_2S_2S_4_2793_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2818_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_Minus_2S_2S_4_2793_out1)
          begin :bnn_N_Mux_2_2_3_4_2819
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2819_out1 = bnn_Minus_2S_2S_4_2793_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2819_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2015_out1 or bnn_Minus_2S_2S_4_2766_out1)
          begin :bnn_N_Mux_2_2_3_4_2820
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2820_out1 = bnn_Minus_2S_2S_4_2766_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2820_out1 = bnn_N_Mux_2_2_3_1_2015_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2821
         assign bnn_Minus_2S_2S_4_2821_out1 = -bnn_N_Mux_2_2_3_1_2049_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_17_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4794_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2824_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2824_in2 = {bnn_Mul_16Sx12S_19S_4_4794_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2824_in2 = {{ 5 {fixed_buffer_17_if_1_dout_wire[11]}}, fixed_buffer_17_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2798_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2824_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2824_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2824_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2798_out1[4]}}, bnn_Add_5Sx4S_6S_1_2798_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2824
         assign bnn_Add_17Sx16S_17S_1_2824_out1 = bnn_Add_17Sx16S_17S_1_2824_in2 + {bnn_Add_17Sx16S_17S_1_2824_in1[15], bnn_Add_17Sx16S_17S_1_2824_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2825
         assign bnn_Add_5Sx4S_6S_1_2825_out1 = {bnn_Add_5Sx4S_6S_1_2800_out1[4], bnn_Add_5Sx4S_6S_1_2800_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2799_out1[1]}}, bnn_N_Mux_2_2_3_4_2799_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2086_out1 or bnn_Minus_2S_2S_4_2801_out1)
          begin :bnn_N_Mux_2_2_3_4_2826
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2826_out1 = bnn_Minus_2S_2S_4_2801_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2826_out1 = bnn_N_Mux_2_2_3_1_2086_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2827
         assign bnn_Add_5Sx4S_6S_1_2827_out1 = {bnn_Add_5Sx4S_6S_1_2803_out1[4], bnn_Add_5Sx4S_6S_1_2803_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2802_out1[1]}}, bnn_N_Mux_2_2_3_4_2802_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2828
         assign bnn_Minus_2S_2S_4_2828_out1 = -bnn_N_Mux_2_2_3_1_2103_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2086_out1 or bnn_Minus_2S_2S_4_2801_out1)
          begin :bnn_N_Mux_2_2_3_4_2829
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2829_out1 = bnn_Minus_2S_2S_4_2801_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2829_out1 = bnn_N_Mux_2_2_3_1_2086_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2830
         assign bnn_Add_5Sx4S_6S_1_2830_out1 = {bnn_Add_4Sx2S_5S_1_2806_out1[4], bnn_Add_4Sx2S_5S_1_2806_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2805_out1[1]}}, bnn_N_Mux_2_2_3_4_2805_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2086_out1 or bnn_Minus_2S_2S_4_2801_out1)
          begin :bnn_N_Mux_2_2_3_4_2832
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2832_out1 = bnn_Minus_2S_2S_4_2801_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2832_out1 = bnn_N_Mux_2_2_3_1_2086_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2833
         assign bnn_Add_4Sx2S_5S_1_2833_out1 = {bnn_Add_4Sx3S_4S_1_2809_out1[3], bnn_Add_4Sx3S_4S_1_2809_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2808_out1[1]}}, bnn_N_Mux_2_2_3_4_2808_out1};

         assign bnn_N_Mux_2_2_3_4_2835_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[23], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2810_out1 or bnn_N_Mux_2_2_3_4_2835_in3)
          begin :bnn_N_Mux_2_2_3_4_2835
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2835_out1 = bnn_Minus_2S_2S_4_2810_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2835_out1 = bnn_N_Mux_2_2_3_4_2835_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2836
         assign bnn_Add_4Sx3S_4S_1_2836_out1 = bnn_Add_4Sx3S_4S_1_2812_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2811_out1[1]}}, bnn_N_Mux_2_2_3_4_2811_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2837
         assign bnn_Minus_2S_2S_4_2837_out1 = -bnn_N_Mux_3_2_6_4_2796_out1_slice;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2810_out1 or bnn_N_Mux_2_2_3_4_2835_in3)
          begin :bnn_N_Mux_2_2_3_4_2838
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2838_out1 = bnn_Minus_2S_2S_4_2810_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2838_out1 = bnn_N_Mux_2_2_3_4_2835_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2839
         assign bnn_Add_4Sx3S_4S_1_2839_out1 = bnn_Add_3Sx3S_4S_1_2815_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2814_out1[1]}}, bnn_N_Mux_2_2_3_4_2814_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2840
         assign bnn_Minus_2S_2S_4_2840_out1 = -bnn_N_Mux_2_4_8_1_2022_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2816_out1 or bnn_N_Mux_3_2_6_4_2768_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2841
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2841_out1 = bnn_Minus_2S_2S_4_2816_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2841_out1 = bnn_N_Mux_3_2_6_4_2768_out1_slice;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2842
         assign bnn_Add_3Sx3S_4S_1_2842_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2818_out1[1]}}, bnn_N_Mux_2_2_3_4_2818_out1} + {bnn_Add_2Sx2S_3S_1_2817_out1[2], bnn_Add_2Sx2S_3S_1_2817_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2844
         assign bnn_Add_2Sx2S_3S_1_2844_out1 = {bnn_N_Mux_2_2_3_4_2820_out1[1], bnn_N_Mux_2_2_3_4_2820_out1} + {bnn_N_Mux_2_2_3_4_2819_out1[1], bnn_N_Mux_2_2_3_4_2819_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_Minus_2S_2S_4_2821_out1)
          begin :bnn_N_Mux_2_2_3_4_2845
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2845_out1 = bnn_Minus_2S_2S_4_2821_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2845_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_Minus_2S_2S_4_2821_out1)
          begin :bnn_N_Mux_2_2_3_4_2846
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2846_out1 = bnn_Minus_2S_2S_4_2821_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2846_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2032_out1 or bnn_Minus_2S_2S_4_2793_out1)
          begin :bnn_N_Mux_2_2_3_4_2847
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2847_out1 = bnn_Minus_2S_2S_4_2793_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2847_out1 = bnn_N_Mux_2_2_3_1_2032_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2848
         assign bnn_Minus_2S_2S_4_2848_out1 = -bnn_N_Mux_2_2_3_1_2066_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_18_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4798_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2851_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2851_in2 = {bnn_Mul_16Sx12S_19S_4_4798_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2851_in2 = {{ 5 {fixed_buffer_18_if_1_dout_wire[11]}}, fixed_buffer_18_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2825_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2851_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2851_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2851_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2825_out1[4]}}, bnn_Add_5Sx4S_6S_1_2825_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2851
         assign bnn_Add_17Sx16S_17S_1_2851_out1 = bnn_Add_17Sx16S_17S_1_2851_in2 + {bnn_Add_17Sx16S_17S_1_2851_in1[15], bnn_Add_17Sx16S_17S_1_2851_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2852
         assign bnn_Add_5Sx4S_6S_1_2852_out1 = {bnn_Add_5Sx4S_6S_1_2827_out1[4], bnn_Add_5Sx4S_6S_1_2827_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2826_out1[1]}}, bnn_N_Mux_2_2_3_4_2826_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2103_out1 or bnn_Minus_2S_2S_4_2828_out1)
          begin :bnn_N_Mux_2_2_3_4_2853
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2853_out1 = bnn_Minus_2S_2S_4_2828_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2853_out1 = bnn_N_Mux_2_2_3_1_2103_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2854
         assign bnn_Add_5Sx4S_6S_1_2854_out1 = {bnn_Add_5Sx4S_6S_1_2830_out1[4], bnn_Add_5Sx4S_6S_1_2830_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2829_out1[1]}}, bnn_N_Mux_2_2_3_4_2829_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2855
         assign bnn_Minus_2S_2S_4_2855_out1 = -bnn_N_Mux_2_2_3_1_2120_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2103_out1 or bnn_Minus_2S_2S_4_2828_out1)
          begin :bnn_N_Mux_2_2_3_4_2856
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2856_out1 = bnn_Minus_2S_2S_4_2828_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2856_out1 = bnn_N_Mux_2_2_3_1_2103_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2857
         assign bnn_Add_5Sx4S_6S_1_2857_out1 = {bnn_Add_4Sx2S_5S_1_2833_out1[4], bnn_Add_4Sx2S_5S_1_2833_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2832_out1[1]}}, bnn_N_Mux_2_2_3_4_2832_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2103_out1 or bnn_Minus_2S_2S_4_2828_out1)
          begin :bnn_N_Mux_2_2_3_4_2859
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2859_out1 = bnn_Minus_2S_2S_4_2828_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2859_out1 = bnn_N_Mux_2_2_3_1_2103_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2860
         assign bnn_Add_4Sx2S_5S_1_2860_out1 = {bnn_Add_4Sx3S_4S_1_2836_out1[3], bnn_Add_4Sx3S_4S_1_2836_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2835_out1[1]}}, bnn_N_Mux_2_2_3_4_2835_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2837_out1 or bnn_N_Mux_3_2_6_4_2796_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_2862
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2862_out1 = bnn_Minus_2S_2S_4_2837_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2862_out1 = bnn_N_Mux_3_2_6_4_2796_out1_slice;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2863
         assign bnn_Add_4Sx3S_4S_1_2863_out1 = bnn_Add_4Sx3S_4S_1_2839_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2838_out1[1]}}, bnn_N_Mux_2_2_3_4_2838_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2864
         assign bnn_Minus_2S_2S_4_2864_out1 = -bnn_N_Mux_2_4_8_1_2039_in3;

         assign bnn_N_Mux_2_2_3_4_2865_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[24], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2840_out1 or bnn_N_Mux_2_2_3_4_2865_in3)
          begin :bnn_N_Mux_2_2_3_4_2865
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2865_out1 = bnn_Minus_2S_2S_4_2840_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2865_out1 = bnn_N_Mux_2_2_3_4_2865_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2866
         assign bnn_Add_4Sx3S_4S_1_2866_out1 = bnn_Add_3Sx3S_4S_1_2842_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2841_out1[1]}}, bnn_N_Mux_2_2_3_4_2841_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2840_out1 or bnn_N_Mux_2_2_3_4_2865_in3)
          begin :bnn_N_Mux_2_2_3_4_2868
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2868_out1 = bnn_Minus_2S_2S_4_2840_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2868_out1 = bnn_N_Mux_2_2_3_4_2865_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2869
         assign bnn_Add_3Sx3S_4S_1_2869_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2845_out1[1]}}, bnn_N_Mux_2_2_3_4_2845_out1} + {bnn_Add_2Sx2S_3S_1_2844_out1[2], bnn_Add_2Sx2S_3S_1_2844_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2871
         assign bnn_Add_2Sx2S_3S_1_2871_out1 = {bnn_N_Mux_2_2_3_4_2847_out1[1], bnn_N_Mux_2_2_3_4_2847_out1} + {bnn_N_Mux_2_2_3_4_2846_out1[1], bnn_N_Mux_2_2_3_4_2846_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_Minus_2S_2S_4_2848_out1)
          begin :bnn_N_Mux_2_2_3_4_2872
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2872_out1 = bnn_Minus_2S_2S_4_2848_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2872_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_Minus_2S_2S_4_2848_out1)
          begin :bnn_N_Mux_2_2_3_4_2873
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2873_out1 = bnn_Minus_2S_2S_4_2848_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2873_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2049_out1 or bnn_Minus_2S_2S_4_2821_out1)
          begin :bnn_N_Mux_2_2_3_4_2874
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2874_out1 = bnn_Minus_2S_2S_4_2821_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2874_out1 = bnn_N_Mux_2_2_3_1_2049_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2875
         assign bnn_Minus_2S_2S_4_2875_out1 = -bnn_N_Mux_2_2_3_1_2083_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_19_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4802_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2878_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2878_in2 = {bnn_Mul_16Sx12S_19S_4_4802_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2878_in2 = {{ 5 {fixed_buffer_19_if_1_dout_wire[11]}}, fixed_buffer_19_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2852_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2878_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2878_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2878_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2852_out1[4]}}, bnn_Add_5Sx4S_6S_1_2852_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2878
         assign bnn_Add_17Sx16S_17S_1_2878_out1 = bnn_Add_17Sx16S_17S_1_2878_in2 + {bnn_Add_17Sx16S_17S_1_2878_in1[15], bnn_Add_17Sx16S_17S_1_2878_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2879
         assign bnn_Add_5Sx4S_6S_1_2879_out1 = {bnn_Add_5Sx4S_6S_1_2854_out1[4], bnn_Add_5Sx4S_6S_1_2854_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2853_out1[1]}}, bnn_N_Mux_2_2_3_4_2853_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2120_out1 or bnn_Minus_2S_2S_4_2855_out1)
          begin :bnn_N_Mux_2_2_3_4_2880
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2880_out1 = bnn_Minus_2S_2S_4_2855_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2880_out1 = bnn_N_Mux_2_2_3_1_2120_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2881
         assign bnn_Add_5Sx4S_6S_1_2881_out1 = {bnn_Add_5Sx4S_6S_1_2857_out1[4], bnn_Add_5Sx4S_6S_1_2857_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2856_out1[1]}}, bnn_N_Mux_2_2_3_4_2856_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2882
         assign bnn_Minus_2S_2S_4_2882_out1 = -bnn_N_Mux_2_2_3_1_2137_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2120_out1 or bnn_Minus_2S_2S_4_2855_out1)
          begin :bnn_N_Mux_2_2_3_4_2883
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2883_out1 = bnn_Minus_2S_2S_4_2855_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2883_out1 = bnn_N_Mux_2_2_3_1_2120_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2884
         assign bnn_Add_5Sx4S_6S_1_2884_out1 = {bnn_Add_4Sx2S_5S_1_2860_out1[4], bnn_Add_4Sx2S_5S_1_2860_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2859_out1[1]}}, bnn_N_Mux_2_2_3_4_2859_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2120_out1 or bnn_Minus_2S_2S_4_2855_out1)
          begin :bnn_N_Mux_2_2_3_4_2886
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2886_out1 = bnn_Minus_2S_2S_4_2855_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2886_out1 = bnn_N_Mux_2_2_3_1_2120_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2887
         assign bnn_Add_4Sx2S_5S_1_2887_out1 = {bnn_Add_4Sx3S_4S_1_2863_out1[3], bnn_Add_4Sx3S_4S_1_2863_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2862_out1[1]}}, bnn_N_Mux_2_2_3_4_2862_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2888
         assign bnn_Minus_2S_2S_4_2888_out1 = -bnn_N_Mux_2_2_3_1_2211_out1;

         assign bnn_N_Mux_2_2_3_4_2889_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[25], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2864_out1 or bnn_N_Mux_2_2_3_4_2889_in3)
          begin :bnn_N_Mux_2_2_3_4_2889
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2889_out1 = bnn_Minus_2S_2S_4_2864_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2889_out1 = bnn_N_Mux_2_2_3_4_2889_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2890
         assign bnn_Add_4Sx3S_4S_1_2890_out1 = bnn_Add_4Sx3S_4S_1_2866_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2865_out1[1]}}, bnn_N_Mux_2_2_3_4_2865_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2891
         assign bnn_Minus_2S_2S_4_2891_out1 = -bnn_N_Mux_2_4_8_1_2056_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2864_out1 or bnn_N_Mux_2_2_3_4_2889_in3)
          begin :bnn_N_Mux_2_2_3_4_2892
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2892_out1 = bnn_Minus_2S_2S_4_2864_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2892_out1 = bnn_N_Mux_2_2_3_4_2889_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2893
         assign bnn_Add_4Sx3S_4S_1_2893_out1 = bnn_Add_3Sx3S_4S_1_2869_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2868_out1[1]}}, bnn_N_Mux_2_2_3_4_2868_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2864_out1 or bnn_N_Mux_2_2_3_4_2889_in3)
          begin :bnn_N_Mux_2_2_3_4_2895
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2895_out1 = bnn_Minus_2S_2S_4_2864_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2895_out1 = bnn_N_Mux_2_2_3_4_2889_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2896
         assign bnn_Add_3Sx3S_4S_1_2896_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2872_out1[1]}}, bnn_N_Mux_2_2_3_4_2872_out1} + {bnn_Add_2Sx2S_3S_1_2871_out1[2], bnn_Add_2Sx2S_3S_1_2871_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2898
         assign bnn_Add_2Sx2S_3S_1_2898_out1 = {bnn_N_Mux_2_2_3_4_2874_out1[1], bnn_N_Mux_2_2_3_4_2874_out1} + {bnn_N_Mux_2_2_3_4_2873_out1[1], bnn_N_Mux_2_2_3_4_2873_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_Minus_2S_2S_4_2875_out1)
          begin :bnn_N_Mux_2_2_3_4_2899
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2899_out1 = bnn_Minus_2S_2S_4_2875_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2899_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_Minus_2S_2S_4_2875_out1)
          begin :bnn_N_Mux_2_2_3_4_2900
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2900_out1 = bnn_Minus_2S_2S_4_2875_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2900_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2066_out1 or bnn_Minus_2S_2S_4_2848_out1)
          begin :bnn_N_Mux_2_2_3_4_2901
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2901_out1 = bnn_Minus_2S_2S_4_2848_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2901_out1 = bnn_N_Mux_2_2_3_1_2066_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2902
         assign bnn_Minus_2S_2S_4_2902_out1 = -bnn_N_Mux_2_2_3_1_2100_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_20_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4806_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2905_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2905_in2 = {bnn_Mul_16Sx12S_19S_4_4806_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2905_in2 = {{ 5 {fixed_buffer_20_if_1_dout_wire[11]}}, fixed_buffer_20_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2879_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2905_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2905_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2905_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2879_out1[4]}}, bnn_Add_5Sx4S_6S_1_2879_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2905
         assign bnn_Add_17Sx16S_17S_1_2905_out1 = bnn_Add_17Sx16S_17S_1_2905_in2 + {bnn_Add_17Sx16S_17S_1_2905_in1[15], bnn_Add_17Sx16S_17S_1_2905_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2906
         assign bnn_Add_5Sx4S_6S_1_2906_out1 = {bnn_Add_5Sx4S_6S_1_2881_out1[4], bnn_Add_5Sx4S_6S_1_2881_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2880_out1[1]}}, bnn_N_Mux_2_2_3_4_2880_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2137_out1 or bnn_Minus_2S_2S_4_2882_out1)
          begin :bnn_N_Mux_2_2_3_4_2907
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2907_out1 = bnn_Minus_2S_2S_4_2882_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2907_out1 = bnn_N_Mux_2_2_3_1_2137_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2908
         assign bnn_Add_5Sx4S_6S_1_2908_out1 = {bnn_Add_5Sx4S_6S_1_2884_out1[4], bnn_Add_5Sx4S_6S_1_2884_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2883_out1[1]}}, bnn_N_Mux_2_2_3_4_2883_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2909
         assign bnn_Minus_2S_2S_4_2909_out1 = -bnn_N_Mux_2_2_3_1_2193_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2137_out1 or bnn_Minus_2S_2S_4_2882_out1)
          begin :bnn_N_Mux_2_2_3_4_2910
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2910_out1 = bnn_Minus_2S_2S_4_2882_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2910_out1 = bnn_N_Mux_2_2_3_1_2137_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2911
         assign bnn_Add_5Sx4S_6S_1_2911_out1 = {bnn_Add_4Sx2S_5S_1_2887_out1[4], bnn_Add_4Sx2S_5S_1_2887_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2886_out1[1]}}, bnn_N_Mux_2_2_3_4_2886_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2912
         assign bnn_Minus_2S_2S_4_2912_out1 = -bnn_N_Mux_2_2_3_1_2024_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2211_out1 or bnn_Minus_2S_2S_4_2888_out1)
          begin :bnn_N_Mux_2_2_3_4_2913
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2913_out1 = bnn_Minus_2S_2S_4_2888_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2913_out1 = bnn_N_Mux_2_2_3_1_2211_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2914
         assign bnn_Add_4Sx2S_5S_1_2914_out1 = {bnn_Add_4Sx3S_4S_1_2890_out1[3], bnn_Add_4Sx3S_4S_1_2890_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2889_out1[1]}}, bnn_N_Mux_2_2_3_4_2889_out1};

         assign bnn_N_Mux_2_2_3_4_2916_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[26], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2891_out1 or bnn_N_Mux_2_2_3_4_2916_in3)
          begin :bnn_N_Mux_2_2_3_4_2916
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2916_out1 = bnn_Minus_2S_2S_4_2891_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2916_out1 = bnn_N_Mux_2_2_3_4_2916_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2917
         assign bnn_Add_4Sx3S_4S_1_2917_out1 = bnn_Add_4Sx3S_4S_1_2893_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2892_out1[1]}}, bnn_N_Mux_2_2_3_4_2892_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2918
         assign bnn_Minus_2S_2S_4_2918_out1 = -bnn_N_Mux_2_4_8_1_2073_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2891_out1 or bnn_N_Mux_2_2_3_4_2916_in3)
          begin :bnn_N_Mux_2_2_3_4_2919
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2919_out1 = bnn_Minus_2S_2S_4_2891_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2919_out1 = bnn_N_Mux_2_2_3_4_2916_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2920
         assign bnn_Add_4Sx3S_4S_1_2920_out1 = bnn_Add_3Sx3S_4S_1_2896_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2895_out1[1]}}, bnn_N_Mux_2_2_3_4_2895_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2891_out1 or bnn_N_Mux_2_2_3_4_2916_in3)
          begin :bnn_N_Mux_2_2_3_4_2922
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2922_out1 = bnn_Minus_2S_2S_4_2891_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2922_out1 = bnn_N_Mux_2_2_3_4_2916_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2923
         assign bnn_Add_3Sx3S_4S_1_2923_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2899_out1[1]}}, bnn_N_Mux_2_2_3_4_2899_out1} + {bnn_Add_2Sx2S_3S_1_2898_out1[2], bnn_Add_2Sx2S_3S_1_2898_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2925
         assign bnn_Add_2Sx2S_3S_1_2925_out1 = {bnn_N_Mux_2_2_3_4_2901_out1[1], bnn_N_Mux_2_2_3_4_2901_out1} + {bnn_N_Mux_2_2_3_4_2900_out1[1], bnn_N_Mux_2_2_3_4_2900_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_Minus_2S_2S_4_2902_out1)
          begin :bnn_N_Mux_2_2_3_4_2926
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2926_out1 = bnn_Minus_2S_2S_4_2902_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2926_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_Minus_2S_2S_4_2902_out1)
          begin :bnn_N_Mux_2_2_3_4_2927
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2927_out1 = bnn_Minus_2S_2S_4_2902_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2927_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2083_out1 or bnn_Minus_2S_2S_4_2875_out1)
          begin :bnn_N_Mux_2_2_3_4_2928
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2928_out1 = bnn_Minus_2S_2S_4_2875_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2928_out1 = bnn_N_Mux_2_2_3_1_2083_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2929
         assign bnn_Minus_2S_2S_1_2929_out1 = -bnn_N_Mux_2_2_3_1_2117_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_21_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4810_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2932_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2932_in2 = {bnn_Mul_16Sx12S_19S_4_4810_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2932_in2 = {{ 5 {fixed_buffer_21_if_1_dout_wire[11]}}, fixed_buffer_21_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2906_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2932_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2932_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2932_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2906_out1[4]}}, bnn_Add_5Sx4S_6S_1_2906_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2932
         assign bnn_Add_17Sx16S_17S_1_2932_out1 = bnn_Add_17Sx16S_17S_1_2932_in2 + {bnn_Add_17Sx16S_17S_1_2932_in1[15], bnn_Add_17Sx16S_17S_1_2932_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2933
         assign bnn_Add_5Sx4S_6S_1_2933_out1 = {bnn_Add_5Sx4S_6S_1_2908_out1[4], bnn_Add_5Sx4S_6S_1_2908_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2907_out1[1]}}, bnn_N_Mux_2_2_3_4_2907_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2193_out1 or bnn_Minus_2S_2S_4_2909_out1)
          begin :bnn_N_Mux_2_2_3_4_2934
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2934_out1 = bnn_Minus_2S_2S_4_2909_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2934_out1 = bnn_N_Mux_2_2_3_1_2193_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2935
         assign bnn_Add_5Sx4S_6S_1_2935_out1 = {bnn_Add_5Sx4S_6S_1_2911_out1[4], bnn_Add_5Sx4S_6S_1_2911_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2910_out1[1]}}, bnn_N_Mux_2_2_3_4_2910_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2936
         assign bnn_Minus_2S_2S_4_2936_out1 = -bnn_N_Mux_2_2_3_1_2041_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2024_out1 or bnn_Minus_2S_2S_4_2912_out1)
          begin :bnn_N_Mux_2_2_3_4_2937
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2937_out1 = bnn_Minus_2S_2S_4_2912_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2937_out1 = bnn_N_Mux_2_2_3_1_2024_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2938
         assign bnn_Add_5Sx4S_6S_1_2938_out1 = {bnn_Add_4Sx2S_5S_1_2914_out1[4], bnn_Add_4Sx2S_5S_1_2914_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2913_out1[1]}}, bnn_N_Mux_2_2_3_4_2913_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2024_out1 or bnn_Minus_2S_2S_4_2912_out1)
          begin :bnn_N_Mux_2_2_3_4_2940
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2940_out1 = bnn_Minus_2S_2S_4_2912_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2940_out1 = bnn_N_Mux_2_2_3_1_2024_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2941
         assign bnn_Add_4Sx2S_5S_1_2941_out1 = {bnn_Add_4Sx3S_4S_1_2917_out1[3], bnn_Add_4Sx3S_4S_1_2917_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2916_out1[1]}}, bnn_N_Mux_2_2_3_4_2916_out1};

         assign bnn_N_Mux_2_2_3_4_2943_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[27], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2918_out1 or bnn_N_Mux_2_2_3_4_2943_in3)
          begin :bnn_N_Mux_2_2_3_4_2943
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2943_out1 = bnn_Minus_2S_2S_4_2918_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2943_out1 = bnn_N_Mux_2_2_3_4_2943_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2944
         assign bnn_Add_4Sx3S_4S_1_2944_out1 = bnn_Add_4Sx3S_4S_1_2920_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2919_out1[1]}}, bnn_N_Mux_2_2_3_4_2919_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2945
         assign bnn_Minus_2S_2S_4_2945_out1 = -bnn_N_Mux_2_4_8_1_2090_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2918_out1 or bnn_N_Mux_2_2_3_4_2943_in3)
          begin :bnn_N_Mux_2_2_3_4_2946
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2946_out1 = bnn_Minus_2S_2S_4_2918_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2946_out1 = bnn_N_Mux_2_2_3_4_2943_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2947
         assign bnn_Add_4Sx3S_4S_1_2947_out1 = bnn_Add_3Sx3S_4S_1_2923_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2922_out1[1]}}, bnn_N_Mux_2_2_3_4_2922_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2918_out1 or bnn_N_Mux_2_2_3_4_2943_in3)
          begin :bnn_N_Mux_2_2_3_4_2949
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2949_out1 = bnn_Minus_2S_2S_4_2918_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2949_out1 = bnn_N_Mux_2_2_3_4_2943_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2950
         assign bnn_Add_3Sx3S_4S_1_2950_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2926_out1[1]}}, bnn_N_Mux_2_2_3_4_2926_out1} + {bnn_Add_2Sx2S_3S_1_2925_out1[2], bnn_Add_2Sx2S_3S_1_2925_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2952
         assign bnn_Add_2Sx2S_3S_1_2952_out1 = {bnn_N_Mux_2_2_3_4_2928_out1[1], bnn_N_Mux_2_2_3_4_2928_out1} + {bnn_N_Mux_2_2_3_4_2927_out1[1], bnn_N_Mux_2_2_3_4_2927_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_Minus_2S_2S_1_2929_out1)
          begin :bnn_N_Mux_2_2_3_4_2953
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2953_out1 = bnn_Minus_2S_2S_1_2929_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2953_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_Minus_2S_2S_1_2929_out1)
          begin :bnn_N_Mux_2_2_3_4_2954
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_4_2954_out1 = bnn_Minus_2S_2S_1_2929_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2954_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2100_out1 or bnn_Minus_2S_2S_4_2902_out1)
          begin :bnn_N_Mux_2_2_3_4_2955
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_4_2955_out1 = bnn_Minus_2S_2S_4_2902_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2955_out1 = bnn_N_Mux_2_2_3_1_2100_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_2956
         assign bnn_Minus_2S_2S_1_2956_out1 = -bnn_N_Mux_2_2_3_1_2134_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_22_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4814_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2957_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2957_in2 = {bnn_Mul_16Sx12S_19S_4_4814_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2957_in2 = {{ 5 {fixed_buffer_22_if_1_dout_wire[11]}}, fixed_buffer_22_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2933_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2957_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2957_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2957_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2933_out1[4]}}, bnn_Add_5Sx4S_6S_1_2933_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2957
         assign bnn_Add_17Sx16S_17S_1_2957_out1 = bnn_Add_17Sx16S_17S_1_2957_in2 + {bnn_Add_17Sx16S_17S_1_2957_in1[15], bnn_Add_17Sx16S_17S_1_2957_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2958
         assign bnn_Add_5Sx4S_6S_1_2958_out1 = {bnn_Add_5Sx4S_6S_1_2935_out1[4], bnn_Add_5Sx4S_6S_1_2935_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2934_out1[1]}}, bnn_N_Mux_2_2_3_4_2934_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2041_out1 or bnn_Minus_2S_2S_4_2936_out1)
          begin :bnn_N_Mux_2_2_3_4_2959
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2959_out1 = bnn_Minus_2S_2S_4_2936_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2959_out1 = bnn_N_Mux_2_2_3_1_2041_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2960
         assign bnn_Add_5Sx4S_6S_1_2960_out1 = {bnn_Add_5Sx4S_6S_1_2938_out1[4], bnn_Add_5Sx4S_6S_1_2938_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2937_out1[1]}}, bnn_N_Mux_2_2_3_4_2937_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2961
         assign bnn_Minus_2S_2S_4_2961_out1 = -bnn_N_Mux_2_2_3_1_2058_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2041_out1 or bnn_Minus_2S_2S_4_2936_out1)
          begin :bnn_N_Mux_2_2_3_4_2962
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2962_out1 = bnn_Minus_2S_2S_4_2936_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2962_out1 = bnn_N_Mux_2_2_3_1_2041_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2963
         assign bnn_Add_5Sx4S_6S_1_2963_out1 = {bnn_Add_4Sx2S_5S_1_2941_out1[4], bnn_Add_4Sx2S_5S_1_2941_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2940_out1[1]}}, bnn_N_Mux_2_2_3_4_2940_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2041_out1 or bnn_Minus_2S_2S_4_2936_out1)
          begin :bnn_N_Mux_2_2_3_4_2965
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2965_out1 = bnn_Minus_2S_2S_4_2936_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2965_out1 = bnn_N_Mux_2_2_3_1_2041_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2966
         assign bnn_Add_4Sx2S_5S_1_2966_out1 = {bnn_Add_4Sx3S_4S_1_2944_out1[3], bnn_Add_4Sx3S_4S_1_2944_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2943_out1[1]}}, bnn_N_Mux_2_2_3_4_2943_out1};

         assign bnn_N_Mux_2_2_3_4_2968_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[28], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2945_out1 or bnn_N_Mux_2_2_3_4_2968_in3)
          begin :bnn_N_Mux_2_2_3_4_2968
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2968_out1 = bnn_Minus_2S_2S_4_2945_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2968_out1 = bnn_N_Mux_2_2_3_4_2968_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2969
         assign bnn_Add_4Sx3S_4S_1_2969_out1 = bnn_Add_4Sx3S_4S_1_2947_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2946_out1[1]}}, bnn_N_Mux_2_2_3_4_2946_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2970
         assign bnn_Minus_2S_2S_4_2970_out1 = -bnn_N_Mux_2_4_8_1_2107_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2945_out1 or bnn_N_Mux_2_2_3_4_2968_in3)
          begin :bnn_N_Mux_2_2_3_4_2971
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2971_out1 = bnn_Minus_2S_2S_4_2945_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2971_out1 = bnn_N_Mux_2_2_3_4_2968_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2972
         assign bnn_Add_4Sx3S_4S_1_2972_out1 = bnn_Add_3Sx3S_4S_1_2950_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2949_out1[1]}}, bnn_N_Mux_2_2_3_4_2949_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2945_out1 or bnn_N_Mux_2_2_3_4_2968_in3)
          begin :bnn_N_Mux_2_2_3_4_2974
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2974_out1 = bnn_Minus_2S_2S_4_2945_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2974_out1 = bnn_N_Mux_2_2_3_4_2968_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2975
         assign bnn_Add_3Sx3S_4S_1_2975_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2953_out1[1]}}, bnn_N_Mux_2_2_3_4_2953_out1} + {bnn_Add_2Sx2S_3S_1_2952_out1[2], bnn_Add_2Sx2S_3S_1_2952_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_2977
         assign bnn_Add_2Sx2S_3S_1_2977_out1 = {bnn_N_Mux_2_2_3_4_2955_out1[1], bnn_N_Mux_2_2_3_4_2955_out1} + {bnn_N_Mux_2_2_3_4_2954_out1[1], bnn_N_Mux_2_2_3_4_2954_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_916 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_Minus_2S_2S_1_2956_out1)
          begin :bnn_N_Mux_2_2_3_4_2978
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_4_2978_out1 = bnn_Minus_2S_2S_1_2956_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2978_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_23_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4818_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2981_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2981_in2 = {bnn_Mul_16Sx12S_19S_4_4818_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2981_in2 = {{ 5 {fixed_buffer_23_if_1_dout_wire[11]}}, fixed_buffer_23_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2958_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_2981_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_2981_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_2981_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2958_out1[4]}}, bnn_Add_5Sx4S_6S_1_2958_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_2981
         assign bnn_Add_17Sx16S_17S_1_2981_out1 = bnn_Add_17Sx16S_17S_1_2981_in2 + {bnn_Add_17Sx16S_17S_1_2981_in1[15], bnn_Add_17Sx16S_17S_1_2981_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2982
         assign bnn_Add_5Sx4S_6S_1_2982_out1 = {bnn_Add_5Sx4S_6S_1_2960_out1[4], bnn_Add_5Sx4S_6S_1_2960_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2959_out1[1]}}, bnn_N_Mux_2_2_3_4_2959_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2058_out1 or bnn_Minus_2S_2S_4_2961_out1)
          begin :bnn_N_Mux_2_2_3_4_2983
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_2983_out1 = bnn_Minus_2S_2S_4_2961_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2983_out1 = bnn_N_Mux_2_2_3_1_2058_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2984
         assign bnn_Add_5Sx4S_6S_1_2984_out1 = {bnn_Add_5Sx4S_6S_1_2963_out1[4], bnn_Add_5Sx4S_6S_1_2963_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2962_out1[1]}}, bnn_N_Mux_2_2_3_4_2962_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2985
         assign bnn_Minus_2S_2S_4_2985_out1 = -bnn_N_Mux_2_2_3_1_2075_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2058_out1 or bnn_Minus_2S_2S_4_2961_out1)
          begin :bnn_N_Mux_2_2_3_4_2986
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_2986_out1 = bnn_Minus_2S_2S_4_2961_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2986_out1 = bnn_N_Mux_2_2_3_1_2058_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_2987
         assign bnn_Add_5Sx4S_6S_1_2987_out1 = {bnn_Add_4Sx2S_5S_1_2966_out1[4], bnn_Add_4Sx2S_5S_1_2966_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2965_out1[1]}}, bnn_N_Mux_2_2_3_4_2965_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2058_out1 or bnn_Minus_2S_2S_4_2961_out1)
          begin :bnn_N_Mux_2_2_3_4_2989
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_2989_out1 = bnn_Minus_2S_2S_4_2961_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2989_out1 = bnn_N_Mux_2_2_3_1_2058_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_2990
         assign bnn_Add_4Sx2S_5S_1_2990_out1 = {bnn_Add_4Sx3S_4S_1_2969_out1[3], bnn_Add_4Sx3S_4S_1_2969_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2968_out1[1]}}, bnn_N_Mux_2_2_3_4_2968_out1};

         assign bnn_N_Mux_2_2_3_4_2992_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[29], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2970_out1 or bnn_N_Mux_2_2_3_4_2992_in3)
          begin :bnn_N_Mux_2_2_3_4_2992
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_2992_out1 = bnn_Minus_2S_2S_4_2970_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2992_out1 = bnn_N_Mux_2_2_3_4_2992_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2993
         assign bnn_Add_4Sx3S_4S_1_2993_out1 = bnn_Add_4Sx3S_4S_1_2972_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2971_out1[1]}}, bnn_N_Mux_2_2_3_4_2971_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_2994
         assign bnn_Minus_2S_2S_4_2994_out1 = -bnn_N_Mux_2_4_8_1_2124_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2970_out1 or bnn_N_Mux_2_2_3_4_2992_in3)
          begin :bnn_N_Mux_2_2_3_4_2995
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_2995_out1 = bnn_Minus_2S_2S_4_2970_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2995_out1 = bnn_N_Mux_2_2_3_4_2992_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_2996
         assign bnn_Add_4Sx3S_4S_1_2996_out1 = bnn_Add_3Sx3S_4S_1_2975_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2974_out1[1]}}, bnn_N_Mux_2_2_3_4_2974_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2970_out1 or bnn_N_Mux_2_2_3_4_2992_in3)
          begin :bnn_N_Mux_2_2_3_4_2998
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_2998_out1 = bnn_Minus_2S_2S_4_2970_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_2998_out1 = bnn_N_Mux_2_2_3_4_2992_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_2999
         assign bnn_Add_3Sx3S_4S_1_2999_out1 = {{ 2 {bnn_N_Mux_2_2_3_4_2978_out1[1]}}, bnn_N_Mux_2_2_3_4_2978_out1} + {bnn_Add_2Sx2S_3S_1_2977_out1[2], bnn_Add_2Sx2S_3S_1_2977_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_907 or bnn_N_Mux_2_2_3_1_2134_out1 or bnn_Minus_2S_2S_1_2956_out1)
          begin :bnn_N_Mux_2_2_3_1_3000
            if (s_reg_907) begin
               bnn_N_Mux_2_2_3_1_3000_out1 = bnn_Minus_2S_2S_1_2956_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3000_out1 = bnn_N_Mux_2_2_3_1_2134_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_908 or bnn_N_Mux_2_2_3_1_2117_out1 or bnn_Minus_2S_2S_1_2929_out1)
          begin :bnn_N_Mux_2_2_3_1_3001
            if (s_reg_908) begin
               bnn_N_Mux_2_2_3_1_3001_out1 = bnn_Minus_2S_2S_1_2929_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3001_out1 = bnn_N_Mux_2_2_3_1_2117_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3002
         assign bnn_Minus_2S_2S_1_3002_out1 = -bnn_N_Mux_3_2_6_1_1783_out1_slice;

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3003
         assign bnn_Minus_2S_2S_1_3003_out1 = -bnn_N_Mux_2_2_3_1_1778_out1;

         // resource: mux_17bx2i
         always @(fixed_buffer_24_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4822_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3005_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3005_in2 = {bnn_Mul_16Sx12S_19S_4_4822_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3005_in2 = {{ 5 {fixed_buffer_24_if_1_dout_wire[11]}}, fixed_buffer_24_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_2982_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3005_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3005_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3005_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_2982_out1[4]}}, bnn_Add_5Sx4S_6S_1_2982_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3005
         assign bnn_Add_17Sx16S_17S_1_3005_out1 = bnn_Add_17Sx16S_17S_1_3005_in2 + {bnn_Add_17Sx16S_17S_1_3005_in1[15], bnn_Add_17Sx16S_17S_1_3005_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3006
         assign bnn_Add_5Sx4S_6S_1_3006_out1 = {bnn_Add_5Sx4S_6S_1_2984_out1[4], bnn_Add_5Sx4S_6S_1_2984_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2983_out1[1]}}, bnn_N_Mux_2_2_3_4_2983_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2075_out1 or bnn_Minus_2S_2S_4_2985_out1)
          begin :bnn_N_Mux_2_2_3_4_3007
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3007_out1 = bnn_Minus_2S_2S_4_2985_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3007_out1 = bnn_N_Mux_2_2_3_1_2075_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3008
         assign bnn_Add_5Sx4S_6S_1_3008_out1 = {bnn_Add_5Sx4S_6S_1_2987_out1[4], bnn_Add_5Sx4S_6S_1_2987_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_2986_out1[1]}}, bnn_N_Mux_2_2_3_4_2986_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3009
         assign bnn_Minus_2S_2S_4_3009_out1 = -bnn_N_Mux_2_2_3_1_2092_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2075_out1 or bnn_Minus_2S_2S_4_2985_out1)
          begin :bnn_N_Mux_2_2_3_4_3010
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3010_out1 = bnn_Minus_2S_2S_4_2985_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3010_out1 = bnn_N_Mux_2_2_3_1_2075_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3011
         assign bnn_Add_5Sx4S_6S_1_3011_out1 = {bnn_Add_4Sx2S_5S_1_2990_out1[4], bnn_Add_4Sx2S_5S_1_2990_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_2989_out1[1]}}, bnn_N_Mux_2_2_3_4_2989_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2075_out1 or bnn_Minus_2S_2S_4_2985_out1)
          begin :bnn_N_Mux_2_2_3_4_3013
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3013_out1 = bnn_Minus_2S_2S_4_2985_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3013_out1 = bnn_N_Mux_2_2_3_1_2075_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_3014
         assign bnn_Add_4Sx2S_5S_1_3014_out1 = {bnn_Add_4Sx3S_4S_1_2993_out1[3], bnn_Add_4Sx3S_4S_1_2993_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_2992_out1[1]}}, bnn_N_Mux_2_2_3_4_2992_out1};

         assign bnn_N_Mux_2_2_3_4_3016_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[30], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_2994_out1 or bnn_N_Mux_2_2_3_4_3016_in3)
          begin :bnn_N_Mux_2_2_3_4_3016
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_3016_out1 = bnn_Minus_2S_2S_4_2994_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3016_out1 = bnn_N_Mux_2_2_3_4_3016_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_3017
         assign bnn_Add_4Sx3S_4S_1_3017_out1 = bnn_Add_4Sx3S_4S_1_2996_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2995_out1[1]}}, bnn_N_Mux_2_2_3_4_2995_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3018
         assign bnn_Minus_2S_2S_4_3018_out1 = -bnn_N_Mux_2_4_8_4_2141_in3;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_2994_out1 or bnn_N_Mux_2_2_3_4_3016_in3)
          begin :bnn_N_Mux_2_2_3_4_3019
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_3019_out1 = bnn_Minus_2S_2S_4_2994_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3019_out1 = bnn_N_Mux_2_2_3_4_3016_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_3020
         assign bnn_Add_4Sx3S_4S_1_3020_out1 = bnn_Add_3Sx3S_4S_1_2999_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_2998_out1[1]}}, bnn_N_Mux_2_2_3_4_2998_out1};

         // resource: bnn_Add_2Sx2S_3S_1  instance: bnn_Add_2Sx2S_3S_1_3022
         assign bnn_Add_2Sx2S_3S_1_3022_out1 = {bnn_N_Mux_2_2_3_1_3001_out1[1], bnn_N_Mux_2_2_3_1_3001_out1} + {bnn_N_Mux_2_2_3_1_3000_out1[1], bnn_N_Mux_2_2_3_1_3000_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_916 or bnn_Minus_2S_2S_1_3002_out1 or bnn_N_Mux_3_2_6_1_1783_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_3023
            if (s_reg_916) begin
               bnn_N_Mux_2_2_3_1_3023_out1 = bnn_Minus_2S_2S_1_3002_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3023_out1 = bnn_N_Mux_3_2_6_1_1783_out1_slice;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3024
         assign bnn_Minus_2S_2S_4_3024_out1 = -bnn_N_Mux_2_2_3_1_1787_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1778_out1 or bnn_Minus_2S_2S_1_3003_out1)
          begin :bnn_N_Mux_2_2_3_4_3025
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3025_out1 = bnn_Minus_2S_2S_1_3003_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3025_out1 = bnn_N_Mux_2_2_3_1_1778_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3026_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[32], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1828_out1 or bnn_N_Mux_2_2_3_1_1831_out1 or bnn_N_Mux_2_2_3_1_1933_out1 or bnn_N_Mux_2_4_8_1_3026_in3)
          begin :bnn_N_Mux_2_4_8_1_3026
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3026_out1 = bnn_N_Mux_2_2_3_1_1828_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3026_out1 = bnn_N_Mux_2_4_8_1_3026_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3026_out1 = bnn_N_Mux_2_2_3_1_1831_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3026_out1 = bnn_N_Mux_2_2_3_1_1933_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1778_out1 or bnn_Minus_2S_2S_1_3003_out1)
          begin :bnn_N_Mux_2_2_3_4_3028
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3028_out1 = bnn_Minus_2S_2S_1_3003_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3028_out1 = bnn_N_Mux_2_2_3_1_1778_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_25_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4826_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3030_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3030_in2 = {bnn_Mul_16Sx12S_19S_4_4826_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3030_in2 = {{ 5 {fixed_buffer_25_if_1_dout_wire[11]}}, fixed_buffer_25_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3006_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3030_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3030_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3030_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3006_out1[4]}}, bnn_Add_5Sx4S_6S_1_3006_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3030
         assign bnn_Add_17Sx16S_17S_1_3030_out1 = bnn_Add_17Sx16S_17S_1_3030_in2 + {bnn_Add_17Sx16S_17S_1_3030_in1[15], bnn_Add_17Sx16S_17S_1_3030_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3031
         assign bnn_Add_5Sx4S_6S_1_3031_out1 = {bnn_Add_5Sx4S_6S_1_3008_out1[4], bnn_Add_5Sx4S_6S_1_3008_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3007_out1[1]}}, bnn_N_Mux_2_2_3_4_3007_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2092_out1 or bnn_Minus_2S_2S_4_3009_out1)
          begin :bnn_N_Mux_2_2_3_4_3032
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3032_out1 = bnn_Minus_2S_2S_4_3009_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3032_out1 = bnn_N_Mux_2_2_3_1_2092_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3033
         assign bnn_Add_5Sx4S_6S_1_3033_out1 = {bnn_Add_5Sx4S_6S_1_3011_out1[4], bnn_Add_5Sx4S_6S_1_3011_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3010_out1[1]}}, bnn_N_Mux_2_2_3_4_3010_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3034
         assign bnn_Minus_2S_2S_4_3034_out1 = -bnn_N_Mux_2_2_3_1_2109_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2092_out1 or bnn_Minus_2S_2S_4_3009_out1)
          begin :bnn_N_Mux_2_2_3_4_3035
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3035_out1 = bnn_Minus_2S_2S_4_3009_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3035_out1 = bnn_N_Mux_2_2_3_1_2092_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3036
         assign bnn_Add_5Sx4S_6S_1_3036_out1 = {bnn_Add_4Sx2S_5S_1_3014_out1[4], bnn_Add_4Sx2S_5S_1_3014_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_3013_out1[1]}}, bnn_N_Mux_2_2_3_4_3013_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2092_out1 or bnn_Minus_2S_2S_4_3009_out1)
          begin :bnn_N_Mux_2_2_3_4_3038
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3038_out1 = bnn_Minus_2S_2S_4_3009_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3038_out1 = bnn_N_Mux_2_2_3_1_2092_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_3039
         assign bnn_Add_4Sx2S_5S_1_3039_out1 = {bnn_Add_4Sx3S_4S_1_3017_out1[3], bnn_Add_4Sx3S_4S_1_3017_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_3016_out1[1]}}, bnn_N_Mux_2_2_3_4_3016_out1};

         assign bnn_N_Mux_2_2_3_4_3041_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[31], 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_939 or bnn_Minus_2S_2S_4_3018_out1 or bnn_N_Mux_2_2_3_4_3041_in3)
          begin :bnn_N_Mux_2_2_3_4_3041
            if (s_reg_939) begin
               bnn_N_Mux_2_2_3_4_3041_out1 = bnn_Minus_2S_2S_4_3018_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3041_out1 = bnn_N_Mux_2_2_3_4_3041_in3;
            end
         end

         // resource: bnn_Add_4Sx3S_4S_1  instance: bnn_Add_4Sx3S_4S_1_3042
         assign bnn_Add_4Sx3S_4S_1_3042_out1 = bnn_Add_4Sx3S_4S_1_3020_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_3019_out1[1]}}, bnn_N_Mux_2_2_3_4_3019_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_924 or bnn_Minus_2S_2S_4_2994_out1 or bnn_N_Mux_2_2_3_4_3016_in3)
          begin :bnn_N_Mux_2_2_3_4_3044
            if (s_reg_924) begin
               bnn_N_Mux_2_2_3_4_3044_out1 = bnn_Minus_2S_2S_4_2994_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3044_out1 = bnn_N_Mux_2_2_3_4_3016_in3;
            end
         end

         // resource: bnn_Add_3Sx3S_4S_1  instance: bnn_Add_3Sx3S_4S_1_3045
         assign bnn_Add_3Sx3S_4S_1_3045_out1 = {{ 2 {bnn_N_Mux_2_2_3_1_3023_out1[1]}}, bnn_N_Mux_2_2_3_1_3023_out1} + {bnn_Add_2Sx2S_3S_1_3022_out1[2], bnn_Add_2Sx2S_3S_1_3022_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1787_out1 or bnn_Minus_2S_2S_4_3024_out1)
          begin :bnn_N_Mux_2_2_3_4_3046
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3046_out1 = bnn_Minus_2S_2S_4_3024_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3046_out1 = bnn_N_Mux_2_2_3_1_1787_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_3047
         assign bnn_Add_5Sx4S_6S_4_3047_out1 = {s_reg_1113[4], s_reg_1113} + {{ 4 {bnn_N_Mux_2_2_3_4_3025_out1[1]}}, bnn_N_Mux_2_2_3_4_3025_out1};

         assign bnn_RightShift_64Sx8S_1S_1_3048_in1 = {s_reg_1032_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3048
         assign bnn_RightShift_64Sx8S_1S_1_3048_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3048_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3026_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3049
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3049_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3049_out1 = bnn_N_Mux_2_4_8_1_3026_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3050_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[33], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1843_out1 or bnn_N_Mux_2_2_3_1_1846_out1 or bnn_N_Mux_2_2_3_1_1944_out1 or bnn_N_Mux_2_4_8_1_3050_in3)
          begin :bnn_N_Mux_2_4_8_1_3050
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3050_out1 = bnn_N_Mux_2_2_3_1_1843_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3050_out1 = bnn_N_Mux_2_4_8_1_3050_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3050_out1 = bnn_N_Mux_2_2_3_1_1846_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3050_out1 = bnn_N_Mux_2_2_3_1_1944_out1;
               end
               
            endcase

         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3051
         assign bnn_Minus_2S_2S_4_3051_out1 = -bnn_N_Mux_2_2_3_1_1792_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1787_out1 or bnn_Minus_2S_2S_4_3024_out1)
          begin :bnn_N_Mux_2_2_3_4_3052
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3052_out1 = bnn_Minus_2S_2S_4_3024_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3052_out1 = bnn_N_Mux_2_2_3_1_1787_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_3053
         assign bnn_Add_5Sx4S_6S_4_3053_out1 = {s_reg_1114[4], s_reg_1114} + {{ 4 {bnn_N_Mux_2_2_3_4_3028_out1[1]}}, bnn_N_Mux_2_2_3_4_3028_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1787_out1 or bnn_Minus_2S_2S_4_3024_out1)
          begin :bnn_N_Mux_2_2_3_4_3055
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3055_out1 = bnn_Minus_2S_2S_4_3024_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3055_out1 = bnn_N_Mux_2_2_3_1_1787_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_26_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4830_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3057_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3057_in2 = {bnn_Mul_16Sx12S_19S_4_4830_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3057_in2 = {{ 5 {fixed_buffer_26_if_1_dout_wire[11]}}, fixed_buffer_26_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3031_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3057_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3057_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3057_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3031_out1[4]}}, bnn_Add_5Sx4S_6S_1_3031_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3057
         assign bnn_Add_17Sx16S_17S_1_3057_out1 = bnn_Add_17Sx16S_17S_1_3057_in2 + {bnn_Add_17Sx16S_17S_1_3057_in1[15], bnn_Add_17Sx16S_17S_1_3057_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3058
         assign bnn_Add_5Sx4S_6S_1_3058_out1 = {bnn_Add_5Sx4S_6S_1_3033_out1[4], bnn_Add_5Sx4S_6S_1_3033_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3032_out1[1]}}, bnn_N_Mux_2_2_3_4_3032_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2109_out1 or bnn_Minus_2S_2S_4_3034_out1)
          begin :bnn_N_Mux_2_2_3_4_3059
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3059_out1 = bnn_Minus_2S_2S_4_3034_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3059_out1 = bnn_N_Mux_2_2_3_1_2109_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3060
         assign bnn_Add_5Sx4S_6S_1_3060_out1 = {bnn_Add_5Sx4S_6S_1_3036_out1[4], bnn_Add_5Sx4S_6S_1_3036_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3035_out1[1]}}, bnn_N_Mux_2_2_3_4_3035_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3061
         assign bnn_Minus_2S_2S_4_3061_out1 = -bnn_N_Mux_2_2_3_1_2126_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2109_out1 or bnn_Minus_2S_2S_4_3034_out1)
          begin :bnn_N_Mux_2_2_3_4_3062
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3062_out1 = bnn_Minus_2S_2S_4_3034_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3062_out1 = bnn_N_Mux_2_2_3_1_2109_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3063
         assign bnn_Add_5Sx4S_6S_1_3063_out1 = {bnn_Add_4Sx2S_5S_1_3039_out1[4], bnn_Add_4Sx2S_5S_1_3039_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_3038_out1[1]}}, bnn_N_Mux_2_2_3_4_3038_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2109_out1 or bnn_Minus_2S_2S_4_3034_out1)
          begin :bnn_N_Mux_2_2_3_4_3065
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3065_out1 = bnn_Minus_2S_2S_4_3034_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3065_out1 = bnn_N_Mux_2_2_3_1_2109_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_3066
         assign bnn_Add_4Sx2S_5S_1_3066_out1 = {bnn_Add_4Sx3S_4S_1_3042_out1[3], bnn_Add_4Sx3S_4S_1_3042_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_3041_out1[1]}}, bnn_N_Mux_2_2_3_4_3041_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_932 or bnn_Minus_2S_2S_4_3018_out1 or bnn_N_Mux_2_2_3_4_3041_in3)
          begin :bnn_N_Mux_2_2_3_4_3068
            if (s_reg_932) begin
               bnn_N_Mux_2_2_3_4_3068_out1 = bnn_Minus_2S_2S_4_3018_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3068_out1 = bnn_N_Mux_2_2_3_4_3041_in3;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_3069
         assign bnn_Add_4Sx2S_4S_1_3069_out1 = bnn_Add_3Sx3S_4S_1_3045_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_3044_out1[1]}}, bnn_N_Mux_2_2_3_4_3044_out1};

         // resource: mux_6bx3i
         always @(s_reg_1130 or bnn_Add_5Sx4S_6S_4_3047_out1[4:0] or bnn_Mod_2Ux32U_7U_4_4450_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_4_3070_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_4_3070_in2 = {s_reg_1130[4], s_reg_1130};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_4_3070_in2 = bnn_Mod_2Ux32U_7U_4_4450_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_4_3070_in2 = {bnn_Add_5Sx4S_6S_4_3047_out1[4], bnn_Add_5Sx4S_6S_4_3047_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1025[1:0] or bnn_N_Mux_2_2_3_4_3046_out1 or bnn_LeftShift_9Ux3U_7U_4_4449_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_4_3070_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_4_3070_in1 = {{ 4 {s_reg_1025[1]}}, s_reg_1025[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_4_3070_in1 = bnn_LeftShift_9Ux3U_7U_4_4449_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_4_3070_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3046_out1[1]}}, bnn_N_Mux_2_2_3_4_3046_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_4  instance: bnn_Add_6Ux6U_6U_4_3070
         assign bnn_Add_6Ux6U_6U_4_3070_out1 = bnn_Add_6Ux6U_6U_4_3070_in2 + bnn_Add_6Ux6U_6U_4_3070_in1;

         assign bnn_N_Mux_2_2_3_1_3071_in3 = {bnn_RightShift_64Sx8S_1S_1_3048_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3049_out1 or bnn_N_Mux_2_2_3_1_3071_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3071
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3071_out1 = bnn_N_Mux_2_2_3_1_3049_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3071_out1 = bnn_N_Mux_2_2_3_1_3071_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3072_in1 = {s_reg_1032_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3072
         assign bnn_RightShift_64Sx8S_1S_1_3072_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3072_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3050_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3073
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3073_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3073_out1 = bnn_N_Mux_2_4_8_1_3050_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3074_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[34], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1854_out1 or bnn_N_Mux_2_2_3_1_1857_out1 or bnn_N_Mux_2_2_3_1_1955_out1 or bnn_N_Mux_2_4_8_1_3074_in3)
          begin :bnn_N_Mux_2_4_8_1_3074
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3074_out1 = bnn_N_Mux_2_2_3_1_1854_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3074_out1 = bnn_N_Mux_2_4_8_1_3074_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3074_out1 = bnn_N_Mux_2_2_3_1_1857_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3074_out1 = bnn_N_Mux_2_2_3_1_1955_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1792_out1 or bnn_Minus_2S_2S_4_3051_out1)
          begin :bnn_N_Mux_2_2_3_4_3075
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3075_out1 = bnn_Minus_2S_2S_4_3051_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3075_out1 = bnn_N_Mux_2_2_3_1_1792_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3076
         assign bnn_Add_5Sx4S_6S_1_3076_out1 = {bnn_Add_5Sx4S_6S_4_3053_out1[4], bnn_Add_5Sx4S_6S_4_3053_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3052_out1[1]}}, bnn_N_Mux_2_2_3_4_3052_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3077
         assign bnn_Minus_2S_2S_4_3077_out1 = -bnn_N_Mux_2_2_3_1_1797_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1792_out1 or bnn_Minus_2S_2S_4_3051_out1)
          begin :bnn_N_Mux_2_2_3_4_3078
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3078_out1 = bnn_Minus_2S_2S_4_3051_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3078_out1 = bnn_N_Mux_2_2_3_1_1792_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3079
         assign bnn_Add_5Sx4S_6S_1_3079_out1 = {s_reg_1115[4], s_reg_1115} + {{ 4 {bnn_N_Mux_2_2_3_4_3055_out1[1]}}, bnn_N_Mux_2_2_3_4_3055_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1792_out1 or bnn_Minus_2S_2S_4_3051_out1)
          begin :bnn_N_Mux_2_2_3_4_3081
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3081_out1 = bnn_Minus_2S_2S_4_3051_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3081_out1 = bnn_N_Mux_2_2_3_1_1792_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_27_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4834_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3083_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3083_in2 = {bnn_Mul_16Sx12S_19S_4_4834_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3083_in2 = {{ 5 {fixed_buffer_27_if_1_dout_wire[11]}}, fixed_buffer_27_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3058_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3083_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3083_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3083_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3058_out1[4]}}, bnn_Add_5Sx4S_6S_1_3058_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3083
         assign bnn_Add_17Sx16S_17S_1_3083_out1 = bnn_Add_17Sx16S_17S_1_3083_in2 + {bnn_Add_17Sx16S_17S_1_3083_in1[15], bnn_Add_17Sx16S_17S_1_3083_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3084
         assign bnn_Add_5Sx4S_6S_1_3084_out1 = {bnn_Add_5Sx4S_6S_1_3060_out1[4], bnn_Add_5Sx4S_6S_1_3060_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3059_out1[1]}}, bnn_N_Mux_2_2_3_4_3059_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2126_out1 or bnn_Minus_2S_2S_4_3061_out1)
          begin :bnn_N_Mux_2_2_3_4_3085
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3085_out1 = bnn_Minus_2S_2S_4_3061_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3085_out1 = bnn_N_Mux_2_2_3_1_2126_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3086
         assign bnn_Add_5Sx4S_6S_1_3086_out1 = {bnn_Add_5Sx4S_6S_1_3063_out1[4], bnn_Add_5Sx4S_6S_1_3063_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3062_out1[1]}}, bnn_N_Mux_2_2_3_4_3062_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3087
         assign bnn_Minus_2S_2S_4_3087_out1 = -bnn_N_Mux_2_2_3_4_2143_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2126_out1 or bnn_Minus_2S_2S_4_3061_out1)
          begin :bnn_N_Mux_2_2_3_4_3088
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3088_out1 = bnn_Minus_2S_2S_4_3061_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3088_out1 = bnn_N_Mux_2_2_3_1_2126_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3089
         assign bnn_Add_5Sx4S_6S_1_3089_out1 = {bnn_Add_4Sx2S_5S_1_3066_out1[4], bnn_Add_4Sx2S_5S_1_3066_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_3065_out1[1]}}, bnn_N_Mux_2_2_3_4_3065_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2126_out1 or bnn_Minus_2S_2S_4_3061_out1)
          begin :bnn_N_Mux_2_2_3_4_3091
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3091_out1 = bnn_Minus_2S_2S_4_3061_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3091_out1 = bnn_N_Mux_2_2_3_1_2126_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_4S_1  instance: bnn_Add_4Sx2S_4S_1_3092
         assign bnn_Add_4Sx2S_4S_1_3092_out1 = bnn_Add_4Sx2S_4S_1_3069_out1 + {{ 2 {bnn_N_Mux_2_2_3_4_3068_out1[1]}}, bnn_N_Mux_2_2_3_4_3068_out1};

         assign bnn_N_Mux_2_2_3_1_3093_in3 = {bnn_RightShift_64Sx8S_1S_1_3072_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3073_out1 or bnn_N_Mux_2_2_3_1_3093_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3093
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3093_out1 = bnn_N_Mux_2_2_3_1_3073_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3093_out1 = bnn_N_Mux_2_2_3_1_3093_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3094_in1 = {s_reg_1032_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3094
         assign bnn_RightShift_64Sx8S_1S_1_3094_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3094_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3074_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3095
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3095_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3095_out1 = bnn_N_Mux_2_4_8_1_3074_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3096_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[35], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1865_out1 or bnn_N_Mux_2_2_3_1_1868_out1 or bnn_N_Mux_2_2_3_1_1966_out1 or bnn_N_Mux_2_4_8_1_3096_in3)
          begin :bnn_N_Mux_2_4_8_1_3096
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3096_out1 = bnn_N_Mux_2_2_3_1_1865_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3096_out1 = bnn_N_Mux_2_4_8_1_3096_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3096_out1 = bnn_N_Mux_2_2_3_1_1868_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3096_out1 = bnn_N_Mux_2_2_3_1_1966_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_32_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4471_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3097_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3097_in2 = {bnn_Mul_16Sx12S_19S_4_4471_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3097_in2 = {{ 5 {fixed_buffer_32_if_1_dout_wire[11]}}, fixed_buffer_32_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_4_3070_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3097_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3097_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3097_in1 = {{ 11 {bnn_Add_6Ux6U_6U_4_3070_out1[4]}}, bnn_Add_6Ux6U_6U_4_3070_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3097
         assign bnn_Add_17Sx16S_17S_1_3097_out1 = bnn_Add_17Sx16S_17S_1_3097_in2 + {bnn_Add_17Sx16S_17S_1_3097_in1[15], bnn_Add_17Sx16S_17S_1_3097_in1};

         // resource: mux_7bx3i
         always @(s_reg_1135 or bnn_Add_5Sx4S_6S_1_3076_out1[4:0] or bnn_Mod_2Ux32U_7U_4_4458_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_7Sx6U_7S_4_3098_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_7Sx6U_7S_4_3098_in2 = {{ 2 {s_reg_1135[4]}}, s_reg_1135};
               end
               
               2'd2: begin
                  bnn_Add_7Sx6U_7S_4_3098_in2 = {1'b0, bnn_Mod_2Ux32U_7U_4_4458_out1[6:1]};
               end
               
               default: begin
                  bnn_Add_7Sx6U_7S_4_3098_in2 = {{ 2 {bnn_Add_5Sx4S_6S_1_3076_out1[4]}}, bnn_Add_5Sx4S_6S_1_3076_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1012[1:0] or bnn_N_Mux_2_2_3_4_3075_out1 or bnn_LeftShift_9Ux3U_7U_4_4457_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_7Sx6U_7S_4_3098_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_7Sx6U_7S_4_3098_in1 = {{ 4 {s_reg_1012[1]}}, s_reg_1012[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_7Sx6U_7S_4_3098_in1 = bnn_LeftShift_9Ux3U_7U_4_4457_out1[6:1];
               end
               
               default: begin
                  bnn_Add_7Sx6U_7S_4_3098_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3075_out1[1]}}, bnn_N_Mux_2_2_3_4_3075_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_7Sx6U_7S_4  instance: bnn_Add_7Sx6U_7S_4_3098
         assign bnn_Add_7Sx6U_7S_4_3098_out1 = bnn_Add_7Sx6U_7S_4_3098_in2 + {1'b0, bnn_Add_7Sx6U_7S_4_3098_in1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1797_out1 or bnn_Minus_2S_2S_4_3077_out1)
          begin :bnn_N_Mux_2_2_3_4_3099
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3099_out1 = bnn_Minus_2S_2S_4_3077_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3099_out1 = bnn_N_Mux_2_2_3_1_1797_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3100
         assign bnn_Add_5Sx4S_6S_1_3100_out1 = {bnn_Add_5Sx4S_6S_1_3079_out1[4], bnn_Add_5Sx4S_6S_1_3079_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3078_out1[1]}}, bnn_N_Mux_2_2_3_4_3078_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3101
         assign bnn_Minus_2S_2S_4_3101_out1 = -bnn_N_Mux_2_2_3_1_1802_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1797_out1 or bnn_Minus_2S_2S_4_3077_out1)
          begin :bnn_N_Mux_2_2_3_4_3102
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3102_out1 = bnn_Minus_2S_2S_4_3077_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3102_out1 = bnn_N_Mux_2_2_3_1_1797_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3103
         assign bnn_Add_5Sx4S_6S_1_3103_out1 = {s_reg_1116[4], s_reg_1116} + {{ 4 {bnn_N_Mux_2_2_3_4_3081_out1[1]}}, bnn_N_Mux_2_2_3_4_3081_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1797_out1 or bnn_Minus_2S_2S_4_3077_out1)
          begin :bnn_N_Mux_2_2_3_4_3105
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3105_out1 = bnn_Minus_2S_2S_4_3077_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3105_out1 = bnn_N_Mux_2_2_3_1_1797_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_28_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4838_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3107_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3107_in2 = {bnn_Mul_16Sx12S_19S_4_4838_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3107_in2 = {{ 5 {fixed_buffer_28_if_1_dout_wire[11]}}, fixed_buffer_28_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3084_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3107_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3107_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3107_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3084_out1[4]}}, bnn_Add_5Sx4S_6S_1_3084_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3107
         assign bnn_Add_17Sx16S_17S_1_3107_out1 = bnn_Add_17Sx16S_17S_1_3107_in2 + {bnn_Add_17Sx16S_17S_1_3107_in1[15], bnn_Add_17Sx16S_17S_1_3107_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3108
         assign bnn_Add_5Sx4S_6S_1_3108_out1 = {bnn_Add_5Sx4S_6S_1_3086_out1[4], bnn_Add_5Sx4S_6S_1_3086_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3085_out1[1]}}, bnn_N_Mux_2_2_3_4_3085_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_4_2143_out1 or bnn_Minus_2S_2S_4_3087_out1)
          begin :bnn_N_Mux_2_2_3_4_3109
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3109_out1 = bnn_Minus_2S_2S_4_3087_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3109_out1 = bnn_N_Mux_2_2_3_4_2143_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3110
         assign bnn_Add_5Sx4S_6S_1_3110_out1 = {bnn_Add_5Sx4S_6S_1_3089_out1[4], bnn_Add_5Sx4S_6S_1_3089_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3088_out1[1]}}, bnn_N_Mux_2_2_3_4_3088_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3111
         assign bnn_Minus_2S_2S_4_3111_out1 = -bnn_N_Mux_3_2_6_1_1785_out1_slice;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_4_2143_out1 or bnn_Minus_2S_2S_4_3087_out1)
          begin :bnn_N_Mux_2_2_3_4_3112
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3112_out1 = bnn_Minus_2S_2S_4_3087_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3112_out1 = bnn_N_Mux_2_2_3_4_2143_out1;
            end
         end

         // resource: bnn_Add_4Sx2S_5S_1  instance: bnn_Add_4Sx2S_5S_1_3113
         assign bnn_Add_4Sx2S_5S_1_3113_out1 = {bnn_Add_4Sx2S_4S_1_3092_out1[3], bnn_Add_4Sx2S_4S_1_3092_out1} + {{ 3 {bnn_N_Mux_2_2_3_4_3091_out1[1]}}, bnn_N_Mux_2_2_3_4_3091_out1};

         assign bnn_N_Mux_2_2_3_1_3114_in3 = {bnn_RightShift_64Sx8S_1S_1_3094_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3095_out1 or bnn_N_Mux_2_2_3_1_3114_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3114
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3114_out1 = bnn_N_Mux_2_2_3_1_3095_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3114_out1 = bnn_N_Mux_2_2_3_1_3114_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3115_in1 = {s_reg_1032_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3115
         assign bnn_RightShift_64Sx8S_1S_1_3115_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3115_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3096_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3116
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3116_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3116_out1 = bnn_N_Mux_2_4_8_1_3096_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3117_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[36], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1876_out1 or bnn_N_Mux_2_2_3_1_1879_out1 or bnn_N_Mux_2_2_3_1_1977_out1 or bnn_N_Mux_2_4_8_1_3117_in3)
          begin :bnn_N_Mux_2_4_8_1_3117
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3117_out1 = bnn_N_Mux_2_2_3_1_1876_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3117_out1 = bnn_N_Mux_2_4_8_1_3117_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3117_out1 = bnn_N_Mux_2_2_3_1_1879_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3117_out1 = bnn_N_Mux_2_2_3_1_1977_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_33_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4433_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3118_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3118_in2 = {bnn_Mul_16Sx12S_19S_4_4433_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3118_in2 = {{ 5 {fixed_buffer_33_if_1_dout_wire[11]}}, fixed_buffer_33_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_7Sx6U_7S_4_3098_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3118_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3118_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3118_in1 = {{ 11 {bnn_Add_7Sx6U_7S_4_3098_out1[4]}}, bnn_Add_7Sx6U_7S_4_3098_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3118
         assign bnn_Add_17Sx16S_17S_1_3118_out1 = bnn_Add_17Sx16S_17S_1_3118_in2 + {bnn_Add_17Sx16S_17S_1_3118_in1[15], bnn_Add_17Sx16S_17S_1_3118_in1};

         // resource: mux_6bx3i
         always @(s_reg_1136 or bnn_Add_5Sx4S_6S_1_3100_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4992_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3119_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3119_in2 = {s_reg_1136[4], s_reg_1136};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3119_in2 = bnn_Mod_6Ux32U_7U_4_4992_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3119_in2 = {bnn_Add_5Sx4S_6S_1_3100_out1[4], bnn_Add_5Sx4S_6S_1_3100_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1030[1:0] or s_reg_1102[6:1] or bnn_N_Mux_2_2_3_4_3099_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3119_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3119_in1 = {{ 4 {s_reg_1030[1]}}, s_reg_1030[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3119_in1 = s_reg_1102[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3119_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3099_out1[1]}}, bnn_N_Mux_2_2_3_4_3099_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3119
         assign bnn_Add_6Ux6U_6U_1_3119_out1 = bnn_Add_6Ux6U_6U_1_3119_in2 + bnn_Add_6Ux6U_6U_1_3119_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1802_out1 or bnn_Minus_2S_2S_4_3101_out1)
          begin :bnn_N_Mux_2_2_3_4_3120
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3120_out1 = bnn_Minus_2S_2S_4_3101_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3120_out1 = bnn_N_Mux_2_2_3_1_1802_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3121
         assign bnn_Add_5Sx4S_6S_1_3121_out1 = {bnn_Add_5Sx4S_6S_1_3103_out1[4], bnn_Add_5Sx4S_6S_1_3103_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3102_out1[1]}}, bnn_N_Mux_2_2_3_4_3102_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3122
         assign bnn_Minus_2S_2S_4_3122_out1 = -bnn_N_Mux_2_2_3_1_1807_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1802_out1 or bnn_Minus_2S_2S_4_3101_out1)
          begin :bnn_N_Mux_2_2_3_4_3123
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3123_out1 = bnn_Minus_2S_2S_4_3101_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3123_out1 = bnn_N_Mux_2_2_3_1_1802_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3124
         assign bnn_Add_5Sx4S_6S_1_3124_out1 = {s_reg_1117[4], s_reg_1117} + {{ 4 {bnn_N_Mux_2_2_3_4_3105_out1[1]}}, bnn_N_Mux_2_2_3_4_3105_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1802_out1 or bnn_Minus_2S_2S_4_3101_out1)
          begin :bnn_N_Mux_2_2_3_4_3126
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3126_out1 = bnn_Minus_2S_2S_4_3101_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3126_out1 = bnn_N_Mux_2_2_3_1_1802_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_29_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4842_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3128_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3128_in2 = {bnn_Mul_16Sx12S_19S_4_4842_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3128_in2 = {{ 5 {fixed_buffer_29_if_1_dout_wire[11]}}, fixed_buffer_29_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3108_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3128_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3128_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3128_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3108_out1[4]}}, bnn_Add_5Sx4S_6S_1_3108_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3128
         assign bnn_Add_17Sx16S_17S_1_3128_out1 = bnn_Add_17Sx16S_17S_1_3128_in2 + {bnn_Add_17Sx16S_17S_1_3128_in1[15], bnn_Add_17Sx16S_17S_1_3128_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3129
         assign bnn_Add_5Sx4S_6S_1_3129_out1 = {bnn_Add_5Sx4S_6S_1_3110_out1[4], bnn_Add_5Sx4S_6S_1_3110_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3109_out1[1]}}, bnn_N_Mux_2_2_3_4_3109_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_4_3111_out1 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_3130
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3130_out1 = bnn_Minus_2S_2S_4_3111_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3130_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3131
         assign bnn_Add_5Sx4S_6S_1_3131_out1 = {bnn_Add_4Sx2S_5S_1_3113_out1[4], bnn_Add_4Sx2S_5S_1_3113_out1} + {{ 4 {bnn_N_Mux_2_2_3_4_3112_out1[1]}}, bnn_N_Mux_2_2_3_4_3112_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3132
         assign bnn_Minus_2S_2S_4_3132_out1 = -bnn_N_Mux_2_2_3_1_1812_out1;

         assign bnn_N_Mux_2_2_3_1_3133_in3 = {bnn_RightShift_64Sx8S_1S_1_3115_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3116_out1 or bnn_N_Mux_2_2_3_1_3133_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3133
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3133_out1 = bnn_N_Mux_2_2_3_1_3116_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3133_out1 = bnn_N_Mux_2_2_3_1_3133_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3134_in1 = {s_reg_1032_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3134
         assign bnn_RightShift_64Sx8S_1S_1_3134_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3134_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3117_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3135
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3135_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3135_out1 = bnn_N_Mux_2_4_8_1_3117_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3136_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[37], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1887_out1 or bnn_N_Mux_2_2_3_1_1890_out1 or bnn_N_Mux_2_2_3_1_1988_out1 or bnn_N_Mux_2_4_8_1_3136_in3)
          begin :bnn_N_Mux_2_4_8_1_3136
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3136_out1 = bnn_N_Mux_2_2_3_1_1887_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3136_out1 = bnn_N_Mux_2_4_8_1_3136_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3136_out1 = bnn_N_Mux_2_2_3_1_1890_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3136_out1 = bnn_N_Mux_2_2_3_1_1988_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_34_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4481_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3137_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3137_in2 = {bnn_Mul_16Sx12S_19S_4_4481_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3137_in2 = {{ 5 {fixed_buffer_34_if_1_dout_wire[11]}}, fixed_buffer_34_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3119_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3137_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3137_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3137_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3119_out1[4]}}, bnn_Add_6Ux6U_6U_1_3119_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3137
         assign bnn_Add_17Sx16S_17S_1_3137_out1 = bnn_Add_17Sx16S_17S_1_3137_in2 + {bnn_Add_17Sx16S_17S_1_3137_in1[15], bnn_Add_17Sx16S_17S_1_3137_in1};

         // resource: mux_6bx3i
         always @(s_reg_1137 or bnn_Add_5Sx4S_6S_1_3121_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4993_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3138_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3138_in2 = {s_reg_1137[4], s_reg_1137};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3138_in2 = bnn_Mod_6Ux32U_7U_4_4993_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3138_in2 = {bnn_Add_5Sx4S_6S_1_3121_out1[4], bnn_Add_5Sx4S_6S_1_3121_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1101[6:1] or s_reg_1108[1:0] or bnn_N_Mux_2_2_3_4_3120_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3138_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3138_in1 = {{ 4 {s_reg_1108[1]}}, s_reg_1108[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3138_in1 = s_reg_1101[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3138_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3120_out1[1]}}, bnn_N_Mux_2_2_3_4_3120_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3138
         assign bnn_Add_6Ux6U_6U_1_3138_out1 = bnn_Add_6Ux6U_6U_1_3138_in2 + bnn_Add_6Ux6U_6U_1_3138_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1807_out1 or bnn_Minus_2S_2S_4_3122_out1)
          begin :bnn_N_Mux_2_2_3_4_3139
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3139_out1 = bnn_Minus_2S_2S_4_3122_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3139_out1 = bnn_N_Mux_2_2_3_1_1807_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3140
         assign bnn_Add_5Sx4S_6S_1_3140_out1 = {bnn_Add_5Sx4S_6S_1_3124_out1[4], bnn_Add_5Sx4S_6S_1_3124_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3123_out1[1]}}, bnn_N_Mux_2_2_3_4_3123_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1807_out1 or bnn_Minus_2S_2S_4_3122_out1)
          begin :bnn_N_Mux_2_2_3_4_3142
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3142_out1 = bnn_Minus_2S_2S_4_3122_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3142_out1 = bnn_N_Mux_2_2_3_1_1807_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3143
         assign bnn_Add_5Sx4S_6S_1_3143_out1 = {s_reg_1118[4], s_reg_1118} + {{ 4 {bnn_N_Mux_2_2_3_4_3126_out1[1]}}, bnn_N_Mux_2_2_3_4_3126_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1807_out1 or bnn_Minus_2S_2S_4_3122_out1)
          begin :bnn_N_Mux_2_2_3_4_3145
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3145_out1 = bnn_Minus_2S_2S_4_3122_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3145_out1 = bnn_N_Mux_2_2_3_1_1807_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_30_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4846_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3146_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3146_in2 = {bnn_Mul_16Sx12S_19S_4_4846_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3146_in2 = {{ 5 {fixed_buffer_30_if_1_dout_wire[11]}}, fixed_buffer_30_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3129_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3146_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3146_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3146_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3129_out1[4]}}, bnn_Add_5Sx4S_6S_1_3129_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3146
         assign bnn_Add_17Sx16S_17S_1_3146_out1 = bnn_Add_17Sx16S_17S_1_3146_in2 + {bnn_Add_17Sx16S_17S_1_3146_in1[15], bnn_Add_17Sx16S_17S_1_3146_in1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3147
         assign bnn_Add_5Sx4S_6S_1_3147_out1 = {bnn_Add_5Sx4S_6S_1_3131_out1[4], bnn_Add_5Sx4S_6S_1_3131_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3130_out1[1]}}, bnn_N_Mux_2_2_3_4_3130_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3148
         assign bnn_Minus_2S_2S_4_3148_out1 = -bnn_N_Mux_2_2_3_1_1817_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1812_out1 or bnn_Minus_2S_2S_4_3132_out1)
          begin :bnn_N_Mux_2_2_3_4_3149
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3149_out1 = bnn_Minus_2S_2S_4_3132_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3149_out1 = bnn_N_Mux_2_2_3_1_1812_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3150
         assign bnn_Minus_2S_2S_1_3150_out1 = -bnn_N_Mux_2_2_3_1_1915_out1;

         assign bnn_N_Mux_2_2_3_1_3151_in3 = {bnn_RightShift_64Sx8S_1S_1_3134_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3135_out1 or bnn_N_Mux_2_2_3_1_3151_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3151
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3151_out1 = bnn_N_Mux_2_2_3_1_3135_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3151_out1 = bnn_N_Mux_2_2_3_1_3151_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3152_in1 = {s_reg_1032_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3152
         assign bnn_RightShift_64Sx8S_1S_1_3152_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3152_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3136_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3153
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3153_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3153_out1 = bnn_N_Mux_2_4_8_1_3136_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3154_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[38], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1898_out1 or bnn_N_Mux_2_2_3_1_1901_out1 or bnn_N_Mux_2_2_3_1_1999_out1 or bnn_N_Mux_2_4_8_1_3154_in3)
          begin :bnn_N_Mux_2_4_8_1_3154
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3154_out1 = bnn_N_Mux_2_2_3_1_1898_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3154_out1 = bnn_N_Mux_2_4_8_1_3154_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3154_out1 = bnn_N_Mux_2_2_3_1_1901_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3154_out1 = bnn_N_Mux_2_2_3_1_1999_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_35_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4491_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3155_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3155_in2 = {bnn_Mul_16Sx12S_19S_4_4491_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3155_in2 = {{ 5 {fixed_buffer_35_if_1_dout_wire[11]}}, fixed_buffer_35_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3138_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3155_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3155_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3155_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3138_out1[4]}}, bnn_Add_6Ux6U_6U_1_3138_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3155
         assign bnn_Add_17Sx16S_17S_1_3155_out1 = bnn_Add_17Sx16S_17S_1_3155_in2 + {bnn_Add_17Sx16S_17S_1_3155_in1[15], bnn_Add_17Sx16S_17S_1_3155_in1};

         // resource: mux_6bx3i
         always @(s_reg_1143 or bnn_Add_5Sx4S_6S_1_3140_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4994_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3156_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3156_in2 = {s_reg_1143[4], s_reg_1143};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3156_in2 = bnn_Mod_6Ux32U_7U_4_4994_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3156_in2 = {bnn_Add_5Sx4S_6S_1_3140_out1[4], bnn_Add_5Sx4S_6S_1_3140_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1099[1:0] or s_reg_886[6:1] or bnn_N_Mux_2_2_3_4_3139_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3156_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3156_in1 = {{ 4 {s_reg_1099[1]}}, s_reg_1099[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3156_in1 = s_reg_886[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3156_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3139_out1[1]}}, bnn_N_Mux_2_2_3_4_3139_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3156
         assign bnn_Add_6Ux6U_6U_1_3156_out1 = bnn_Add_6Ux6U_6U_1_3156_in2 + bnn_Add_6Ux6U_6U_1_3156_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1812_out1 or bnn_Minus_2S_2S_4_3132_out1)
          begin :bnn_N_Mux_2_2_3_4_3157
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3157_out1 = bnn_Minus_2S_2S_4_3132_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3157_out1 = bnn_N_Mux_2_2_3_1_1812_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3158
         assign bnn_Add_5Sx4S_6S_1_3158_out1 = {bnn_Add_5Sx4S_6S_1_3143_out1[4], bnn_Add_5Sx4S_6S_1_3143_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3142_out1[1]}}, bnn_N_Mux_2_2_3_4_3142_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1812_out1 or bnn_Minus_2S_2S_4_3132_out1)
          begin :bnn_N_Mux_2_2_3_4_3160
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3160_out1 = bnn_Minus_2S_2S_4_3132_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3160_out1 = bnn_N_Mux_2_2_3_1_1812_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3161
         assign bnn_Add_5Sx4S_6S_1_3161_out1 = {s_reg_1119[4], s_reg_1119} + {{ 4 {bnn_N_Mux_2_2_3_4_3145_out1[1]}}, bnn_N_Mux_2_2_3_4_3145_out1};

         // resource: mux_17bx2i
         always @(fixed_buffer_31_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4430_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3162_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3162_in2 = {bnn_Mul_16Sx12S_19S_4_4430_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3162_in2 = {{ 5 {fixed_buffer_31_if_1_dout_wire[11]}}, fixed_buffer_31_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_5Sx4S_6S_1_3147_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3162_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3162_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3162_in1 = {{ 11 {bnn_Add_5Sx4S_6S_1_3147_out1[4]}}, bnn_Add_5Sx4S_6S_1_3147_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3162
         assign bnn_Add_17Sx16S_17S_1_3162_out1 = bnn_Add_17Sx16S_17S_1_3162_in2 + {bnn_Add_17Sx16S_17S_1_3162_in1[15], bnn_Add_17Sx16S_17S_1_3162_in1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3163
         assign bnn_Minus_2S_2S_4_3163_out1 = -bnn_N_Mux_2_2_3_1_2149_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1817_out1 or bnn_Minus_2S_2S_4_3148_out1)
          begin :bnn_N_Mux_2_2_3_4_3164
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3164_out1 = bnn_Minus_2S_2S_4_3148_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3164_out1 = bnn_N_Mux_2_2_3_1_1817_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3165
         assign bnn_Add_5Sx4S_6S_1_3165_out1 = {s_reg_1120[4], s_reg_1120} + {{ 4 {bnn_N_Mux_2_2_3_4_3149_out1[1]}}, bnn_N_Mux_2_2_3_4_3149_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3166
         assign bnn_Minus_2S_2S_1_3166_out1 = -bnn_N_Mux_2_2_3_1_1822_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1915_out1 or bnn_Minus_2S_2S_1_3150_out1)
          begin :bnn_N_Mux_2_2_3_1_3167
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3167_out1 = bnn_Minus_2S_2S_1_3150_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3167_out1 = bnn_N_Mux_2_2_3_1_1915_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3168_in3 = {bnn_RightShift_64Sx8S_1S_1_3152_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3153_out1 or bnn_N_Mux_2_2_3_1_3168_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3168
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3168_out1 = bnn_N_Mux_2_2_3_1_3153_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3168_out1 = bnn_N_Mux_2_2_3_1_3168_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3169_in1 = {s_reg_1032_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3169
         assign bnn_RightShift_64Sx8S_1S_1_3169_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3169_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3154_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3170
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3170_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3170_out1 = bnn_N_Mux_2_4_8_1_3154_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3171_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[39], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1909_out1 or bnn_N_Mux_2_2_3_1_1912_out1 or bnn_N_Mux_2_2_3_1_2010_out1 or bnn_N_Mux_2_4_8_4_3171_in3)
          begin :bnn_N_Mux_2_4_8_4_3171
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3171_out1 = bnn_N_Mux_2_2_3_1_1909_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3171_out1 = bnn_N_Mux_2_4_8_4_3171_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3171_out1 = bnn_N_Mux_2_2_3_1_1912_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3171_out1 = bnn_N_Mux_2_2_3_1_2010_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2173_out1 or bnn_N_Mux_2_2_3_1_2176_out1 or bnn_N_Mux_2_2_3_1_2208_out1 or bnn_N_Mux_2_4_8_4_3171_in3)
          begin :bnn_N_Mux_2_4_8_1_3172
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3172_out1 = bnn_N_Mux_2_2_3_1_2173_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3172_out1 = bnn_N_Mux_2_4_8_4_3171_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3172_out1 = bnn_N_Mux_2_2_3_1_2176_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3172_out1 = bnn_N_Mux_2_2_3_1_2208_out1;
               end
               
            endcase

         end

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3173
         assign bnn_RightShift_64Sx8S_1S_1_3173_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_Sub_8Sx2S_8S_4_1600_out1[5:0];

         // resource: mux_17bx2i
         always @(fixed_buffer_36_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4501_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3174_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3174_in2 = {bnn_Mul_16Sx12S_19S_4_4501_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3174_in2 = {{ 5 {fixed_buffer_36_if_1_dout_wire[11]}}, fixed_buffer_36_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3156_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3174_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3174_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3174_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3156_out1[4]}}, bnn_Add_6Ux6U_6U_1_3156_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3174
         assign bnn_Add_17Sx16S_17S_1_3174_out1 = bnn_Add_17Sx16S_17S_1_3174_in2 + {bnn_Add_17Sx16S_17S_1_3174_in1[15], bnn_Add_17Sx16S_17S_1_3174_in1};

         // resource: mux_6bx3i
         always @(s_reg_1035 or bnn_Add_5Sx4S_6S_1_3158_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4995_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3175_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3175_in2 = {s_reg_1035[4], s_reg_1035};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3175_in2 = bnn_Mod_6Ux32U_7U_4_4995_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3175_in2 = {bnn_Add_5Sx4S_6S_1_3158_out1[4], bnn_Add_5Sx4S_6S_1_3158_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1093[6:1] or s_reg_1109[1:0] or bnn_N_Mux_2_2_3_4_3157_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3175_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3175_in1 = {{ 4 {s_reg_1109[1]}}, s_reg_1109[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3175_in1 = s_reg_1093[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3175_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3157_out1[1]}}, bnn_N_Mux_2_2_3_4_3157_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3175
         assign bnn_Add_6Ux6U_6U_1_3175_out1 = bnn_Add_6Ux6U_6U_1_3175_in2 + bnn_Add_6Ux6U_6U_1_3175_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1817_out1 or bnn_Minus_2S_2S_4_3148_out1)
          begin :bnn_N_Mux_2_2_3_4_3176
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3176_out1 = bnn_Minus_2S_2S_4_3148_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3176_out1 = bnn_N_Mux_2_2_3_1_1817_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3177
         assign bnn_Add_5Sx4S_6S_1_3177_out1 = {bnn_Add_5Sx4S_6S_1_3161_out1[4], bnn_Add_5Sx4S_6S_1_3161_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3160_out1[1]}}, bnn_N_Mux_2_2_3_4_3160_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2149_out1 or bnn_Minus_2S_2S_4_3163_out1)
          begin :bnn_N_Mux_2_2_3_4_3179
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3179_out1 = bnn_Minus_2S_2S_4_3163_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3179_out1 = bnn_N_Mux_2_2_3_1_2149_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3180
         assign bnn_Add_5Sx4S_6S_1_3180_out1 = {bnn_Add_5Sx4S_6S_1_3165_out1[4], bnn_Add_5Sx4S_6S_1_3165_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3164_out1[1]}}, bnn_N_Mux_2_2_3_4_3164_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3181
         assign bnn_Minus_2S_2S_1_3181_out1 = -bnn_N_Mux_2_2_3_1_1837_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1822_out1 or bnn_Minus_2S_2S_1_3166_out1)
          begin :bnn_N_Mux_2_2_3_1_3182
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3182_out1 = bnn_Minus_2S_2S_1_3166_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3182_out1 = bnn_N_Mux_2_2_3_1_1822_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3183
         assign bnn_Add_5Sx4S_6S_1_3183_out1 = {s_reg_1121[4], s_reg_1121} + {{ 4 {bnn_N_Mux_2_2_3_1_3167_out1[1]}}, bnn_N_Mux_2_2_3_1_3167_out1};

         assign bnn_N_Mux_2_2_3_1_3184_in3 = {bnn_RightShift_64Sx8S_1S_1_3169_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3170_out1 or bnn_N_Mux_2_2_3_1_3184_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_1_3184
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3184_out1 = bnn_N_Mux_2_2_3_1_3170_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3184_out1 = bnn_N_Mux_2_2_3_1_3184_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3185_in1 = {s_reg_1032_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3185
         assign bnn_RightShift_64Sx8S_1S_4_3185_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3185_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3171_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_4_3186
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_4_3186_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3186_out1 = bnn_N_Mux_2_4_8_4_3171_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3187_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[40], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2161_out1 or bnn_N_Mux_2_2_3_1_2164_out1 or bnn_N_Mux_2_2_3_1_2190_out1 or bnn_N_Mux_2_4_8_1_3187_in3)
          begin :bnn_N_Mux_2_4_8_1_3187
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3187_out1 = bnn_N_Mux_2_2_3_1_2161_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3187_out1 = bnn_N_Mux_2_4_8_1_3187_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3187_out1 = bnn_N_Mux_2_2_3_1_2164_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3187_out1 = bnn_N_Mux_2_2_3_1_2190_out1;
               end
               
            endcase

         end

         assign bnn_RightShift_64Sx8S_1S_1_3188_in1 = {s_reg_1107[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3188
         assign bnn_RightShift_64Sx8S_1S_1_3188_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3188_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3172_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3189
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3189_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3189_out1 = bnn_N_Mux_2_4_8_1_3172_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_1_3190_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_3173_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_3190_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_3190
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_3190_out1_slice = bnn_N_Mux_3_2_6_1_3190_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_3190_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1930_out1 or bnn_N_Mux_2_2_3_1_1933_out1 or bnn_N_Mux_2_2_3_1_2021_out1 or bnn_N_Mux_2_4_8_1_3187_in3)
          begin :bnn_N_Mux_2_4_8_1_3191
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3191_out1 = bnn_N_Mux_2_2_3_1_1930_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3191_out1 = bnn_N_Mux_2_4_8_1_3187_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3191_out1 = bnn_N_Mux_2_2_3_1_1933_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3191_out1 = bnn_N_Mux_2_2_3_1_2021_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_37_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4511_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3192_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3192_in2 = {bnn_Mul_16Sx12S_19S_4_4511_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3192_in2 = {{ 5 {fixed_buffer_37_if_1_dout_wire[11]}}, fixed_buffer_37_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3175_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3192_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3192_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3192_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3175_out1[4]}}, bnn_Add_6Ux6U_6U_1_3175_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3192
         assign bnn_Add_17Sx16S_17S_1_3192_out1 = bnn_Add_17Sx16S_17S_1_3192_in2 + {bnn_Add_17Sx16S_17S_1_3192_in1[15], bnn_Add_17Sx16S_17S_1_3192_in1};

         // resource: mux_6bx3i
         always @(s_reg_1036 or bnn_Add_5Sx4S_6S_1_3177_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4996_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3193_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3193_in2 = {s_reg_1036[4], s_reg_1036};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3193_in2 = bnn_Mod_6Ux32U_7U_4_4996_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3193_in2 = {bnn_Add_5Sx4S_6S_1_3177_out1[4], bnn_Add_5Sx4S_6S_1_3177_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1097[6:1] or s_reg_1110[1:0] or bnn_N_Mux_2_2_3_4_3176_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3193_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3193_in1 = {{ 4 {s_reg_1110[1]}}, s_reg_1110[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3193_in1 = s_reg_1097[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3193_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3176_out1[1]}}, bnn_N_Mux_2_2_3_4_3176_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3193
         assign bnn_Add_6Ux6U_6U_1_3193_out1 = bnn_Add_6Ux6U_6U_1_3193_in2 + bnn_Add_6Ux6U_6U_1_3193_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1822_out1 or bnn_Minus_2S_2S_1_3166_out1)
          begin :bnn_N_Mux_2_2_3_1_3195
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3195_out1 = bnn_Minus_2S_2S_1_3166_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3195_out1 = bnn_N_Mux_2_2_3_1_1822_out1;
            end
         end

         // resource: mux_6bx3i
         always @(s_reg_1039 or bnn_Add_5Sx4S_6S_1_3180_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4997_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3197_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3197_in2 = {s_reg_1039[4], s_reg_1039};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3197_in2 = bnn_Mod_6Ux32U_7U_4_4997_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3197_in2 = {bnn_Add_5Sx4S_6S_1_3180_out1[4], bnn_Add_5Sx4S_6S_1_3180_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1095[6:1] or s_reg_1113[1:0] or bnn_N_Mux_2_2_3_4_3179_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3197_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3197_in1 = {{ 4 {s_reg_1113[1]}}, s_reg_1113[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3197_in1 = s_reg_1095[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3197_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3179_out1[1]}}, bnn_N_Mux_2_2_3_4_3179_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3197
         assign bnn_Add_6Ux6U_6U_1_3197_out1 = bnn_Add_6Ux6U_6U_1_3197_in2 + bnn_Add_6Ux6U_6U_1_3197_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1837_out1 or bnn_Minus_2S_2S_1_3181_out1)
          begin :bnn_N_Mux_2_2_3_4_3198
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3198_out1 = bnn_Minus_2S_2S_1_3181_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3198_out1 = bnn_N_Mux_2_2_3_1_1837_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3183_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5019_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3199_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3199_in2 = bnn_Mod_6Ux32U_7U_4_5019_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3199_in2 = {bnn_Add_5Sx4S_6S_1_3183_out1[4], bnn_Add_5Sx4S_6S_1_3183_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1163[6:1] or bnn_N_Mux_2_2_3_1_3182_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3199_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3199_in1 = s_reg_1163[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3199_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3182_out1[1]}}, bnn_N_Mux_2_2_3_1_3182_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3199
         assign bnn_Add_6Ux6U_6U_1_3199_out1 = bnn_Add_6Ux6U_6U_1_3199_in2 + bnn_Add_6Ux6U_6U_1_3199_in1;

         assign bnn_N_Mux_2_2_3_4_3200_in3 = {bnn_RightShift_64Sx8S_1S_4_3185_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_2_3_4_3186_out1 or bnn_N_Mux_2_2_3_4_3200_in3 or s_reg_1042_stage1)
          begin :bnn_N_Mux_2_2_3_4_3200
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_4_3200_out1 = bnn_N_Mux_2_2_3_4_3186_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3200_out1 = bnn_N_Mux_2_2_3_4_3200_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3187_out1 or s_reg_1056_stage1)
          begin :bnn_N_Mux_2_2_3_1_3201
            if (s_reg_1056_stage1) begin
               bnn_N_Mux_2_2_3_1_3201_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3201_out1 = bnn_N_Mux_2_4_8_1_3187_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_1_3202_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_3188_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_1_3202_in2[1:0])
          begin :bnn_N_Mux_3_2_6_1_3202
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_1_3202_out1_slice = bnn_N_Mux_3_2_6_1_3202_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_3202_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3189_out1 or bnn_N_Mux_3_2_6_1_3190_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_3203
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3203_out1 = bnn_N_Mux_2_2_3_1_3189_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3203_out1 = bnn_N_Mux_3_2_6_1_3190_out1_slice;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3204_in1 = {s_reg_1041_stage1_slice[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3204
         assign bnn_RightShift_64Sx8S_1S_1_3204_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3204_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3191_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3205
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3205_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3205_out1 = bnn_N_Mux_2_4_8_1_3191_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3206_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[41], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1941_out1 or bnn_N_Mux_2_2_3_1_1944_out1 or bnn_N_Mux_2_2_3_1_2038_out1 or bnn_N_Mux_2_4_8_1_3206_in3)
          begin :bnn_N_Mux_2_4_8_1_3206
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3206_out1 = bnn_N_Mux_2_2_3_1_1941_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3206_out1 = bnn_N_Mux_2_4_8_1_3206_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3206_out1 = bnn_N_Mux_2_2_3_1_1944_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3206_out1 = bnn_N_Mux_2_2_3_1_2038_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_38_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4521_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3207_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3207_in2 = {bnn_Mul_16Sx12S_19S_4_4521_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3207_in2 = {{ 5 {fixed_buffer_38_if_1_dout_wire[11]}}, fixed_buffer_38_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3193_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3207_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3207_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3207_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3193_out1[4]}}, bnn_Add_6Ux6U_6U_1_3193_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3207
         assign bnn_Add_17Sx16S_17S_1_3207_out1 = bnn_Add_17Sx16S_17S_1_3207_in2 + {bnn_Add_17Sx16S_17S_1_3207_in1[15], bnn_Add_17Sx16S_17S_1_3207_in1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3208
         assign bnn_Minus_2S_2S_1_3208_out1 = -bnn_N_Mux_2_2_3_1_1848_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1837_out1 or bnn_Minus_2S_2S_1_3181_out1)
          begin :bnn_N_Mux_2_2_3_1_3209
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3209_out1 = bnn_Minus_2S_2S_1_3181_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3209_out1 = bnn_N_Mux_2_2_3_1_1837_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3210
         assign bnn_Add_5Sx4S_6S_1_3210_out1 = {s_reg_1122[4], s_reg_1122} + {{ 4 {bnn_N_Mux_2_2_3_1_3195_out1[1]}}, bnn_N_Mux_2_2_3_1_3195_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1837_out1 or bnn_Minus_2S_2S_1_3181_out1)
          begin :bnn_N_Mux_2_2_3_1_3212
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3212_out1 = bnn_Minus_2S_2S_1_3181_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3212_out1 = bnn_N_Mux_2_2_3_1_1837_out1;
            end
         end

         // resource: mux_6bx3i
         always @(s_reg_1043 or bnn_Add_6Ux6U_6U_1_3199_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4988_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3214_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3214_in2 = {s_reg_1043[4], s_reg_1043};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3214_in2 = bnn_Mod_6Ux32U_7U_4_4988_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3214_in2 = {bnn_Add_6Ux6U_6U_1_3199_out1[4], bnn_Add_6Ux6U_6U_1_3199_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1107[6:1] or s_reg_1114[1:0] or bnn_N_Mux_2_2_3_4_3198_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3214_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3214_in1 = {{ 4 {s_reg_1114[1]}}, s_reg_1114[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3214_in1 = s_reg_1107[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3214_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3198_out1[1]}}, bnn_N_Mux_2_2_3_4_3198_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3214
         assign bnn_Add_6Ux6U_6U_1_3214_out1 = bnn_Add_6Ux6U_6U_1_3214_in2 + bnn_Add_6Ux6U_6U_1_3214_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_2_3_1_3201_out1 or s_reg_1042_stage1 or bnn_N_Mux_3_2_6_1_3202_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_3215
            if (s_reg_1042_stage1) begin
               bnn_N_Mux_2_2_3_1_3215_out1 = bnn_N_Mux_2_2_3_1_3201_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3215_out1 = bnn_N_Mux_3_2_6_1_3202_out1_slice;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3216_in3 = {bnn_RightShift_64Sx8S_1S_1_3204_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3205_out1 or bnn_N_Mux_2_2_3_1_3216_in3)
          begin :bnn_N_Mux_2_2_3_1_3216
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3216_out1 = bnn_N_Mux_2_2_3_1_3205_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3216_out1 = bnn_N_Mux_2_2_3_1_3216_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3217_in1 = {s_reg_1041_stage1_slice[4:0], 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3217
         assign bnn_RightShift_64Sx8S_1S_1_3217_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3217_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3206_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3218
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3218_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3218_out1 = bnn_N_Mux_2_4_8_1_3206_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3219_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[42], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1952_out1 or bnn_N_Mux_2_2_3_1_1955_out1 or bnn_N_Mux_2_2_3_1_2055_out1 or bnn_N_Mux_2_4_8_1_3219_in3)
          begin :bnn_N_Mux_2_4_8_1_3219
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3219_out1 = bnn_N_Mux_2_2_3_1_1952_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3219_out1 = bnn_N_Mux_2_4_8_1_3219_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3219_out1 = bnn_N_Mux_2_2_3_1_1955_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3219_out1 = bnn_N_Mux_2_2_3_1_2055_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_39_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4531_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3220_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3220_in2 = {bnn_Mul_16Sx12S_19S_4_4531_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3220_in2 = {{ 5 {fixed_buffer_39_if_1_dout_wire[11]}}, fixed_buffer_39_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3197_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3220_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3220_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3220_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3197_out1[4]}}, bnn_Add_6Ux6U_6U_1_3197_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3220
         assign bnn_Add_17Sx16S_17S_1_3220_out1 = bnn_Add_17Sx16S_17S_1_3220_in2 + {bnn_Add_17Sx16S_17S_1_3220_in1[15], bnn_Add_17Sx16S_17S_1_3220_in1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1848_out1 or bnn_Minus_2S_2S_1_3208_out1)
          begin :bnn_N_Mux_2_2_3_4_3221
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3221_out1 = bnn_Minus_2S_2S_1_3208_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3221_out1 = bnn_N_Mux_2_2_3_1_1848_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3222
         assign bnn_Add_5Sx4S_6S_1_3222_out1 = {bnn_Add_5Sx4S_6S_1_3210_out1[4], bnn_Add_5Sx4S_6S_1_3210_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3209_out1[1]}}, bnn_N_Mux_2_2_3_1_3209_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3223
         assign bnn_Minus_2S_2S_1_3223_out1 = -bnn_N_Mux_2_2_3_1_1859_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1848_out1 or bnn_Minus_2S_2S_1_3208_out1)
          begin :bnn_N_Mux_2_2_3_1_3224
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3224_out1 = bnn_Minus_2S_2S_1_3208_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3224_out1 = bnn_N_Mux_2_2_3_1_1848_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3225
         assign bnn_Add_5Sx4S_6S_1_3225_out1 = {s_reg_1123[4], s_reg_1123} + {{ 4 {bnn_N_Mux_2_2_3_1_3212_out1[1]}}, bnn_N_Mux_2_2_3_1_3212_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1848_out1 or bnn_Minus_2S_2S_1_3208_out1)
          begin :bnn_N_Mux_2_2_3_1_3227
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3227_out1 = bnn_Minus_2S_2S_1_3208_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3227_out1 = bnn_N_Mux_2_2_3_1_1848_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3229_in3 = {bnn_RightShift_64Sx8S_1S_1_3217_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3218_out1 or bnn_N_Mux_2_2_3_1_3229_in3)
          begin :bnn_N_Mux_2_2_3_1_3229
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3229_out1 = bnn_N_Mux_2_2_3_1_3218_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3229_out1 = bnn_N_Mux_2_2_3_1_3229_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3230_in1 = {s_reg_1041_stage1_slice[4:0], 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3230
         assign bnn_RightShift_64Sx8S_1S_1_3230_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3230_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3219_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3231
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3231_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3231_out1 = bnn_N_Mux_2_4_8_1_3219_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3232_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[43], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1963_out1 or bnn_N_Mux_2_2_3_1_1966_out1 or bnn_N_Mux_2_2_3_1_2072_out1 or bnn_N_Mux_2_4_8_1_3232_in3)
          begin :bnn_N_Mux_2_4_8_1_3232
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3232_out1 = bnn_N_Mux_2_2_3_1_1963_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3232_out1 = bnn_N_Mux_2_4_8_1_3232_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3232_out1 = bnn_N_Mux_2_2_3_1_1966_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3232_out1 = bnn_N_Mux_2_2_3_1_2072_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_40_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4541_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3233_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3233_in2 = {bnn_Mul_16Sx12S_19S_4_4541_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3233_in2 = {{ 5 {fixed_buffer_40_if_1_dout_wire[11]}}, fixed_buffer_40_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3214_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3233_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3233_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3233_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3214_out1[4]}}, bnn_Add_6Ux6U_6U_1_3214_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3233
         assign bnn_Add_17Sx16S_17S_1_3233_out1 = bnn_Add_17Sx16S_17S_1_3233_in2 + {bnn_Add_17Sx16S_17S_1_3233_in1[15], bnn_Add_17Sx16S_17S_1_3233_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3222_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5013_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3234_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3234_in2 = bnn_Mod_6Ux32U_7U_4_5013_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3234_in2 = {bnn_Add_5Sx4S_6S_1_3222_out1[4], bnn_Add_5Sx4S_6S_1_3222_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1103[6:1] or bnn_N_Mux_2_2_3_4_3221_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3234_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3234_in1 = s_reg_1103[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3234_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3221_out1[1]}}, bnn_N_Mux_2_2_3_4_3221_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3234
         assign bnn_Add_6Ux6U_6U_1_3234_out1 = bnn_Add_6Ux6U_6U_1_3234_in2 + bnn_Add_6Ux6U_6U_1_3234_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1859_out1 or bnn_Minus_2S_2S_1_3223_out1)
          begin :bnn_N_Mux_2_2_3_4_3235
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3235_out1 = bnn_Minus_2S_2S_1_3223_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3235_out1 = bnn_N_Mux_2_2_3_1_1859_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3236
         assign bnn_Add_5Sx4S_6S_1_3236_out1 = {bnn_Add_5Sx4S_6S_1_3225_out1[4], bnn_Add_5Sx4S_6S_1_3225_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3224_out1[1]}}, bnn_N_Mux_2_2_3_1_3224_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3237
         assign bnn_Minus_2S_2S_1_3237_out1 = -bnn_N_Mux_2_2_3_1_1870_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1859_out1 or bnn_Minus_2S_2S_1_3223_out1)
          begin :bnn_N_Mux_2_2_3_1_3238
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3238_out1 = bnn_Minus_2S_2S_1_3223_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3238_out1 = bnn_N_Mux_2_2_3_1_1859_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3239
         assign bnn_Add_5Sx4S_6S_1_3239_out1 = {s_reg_1124[4], s_reg_1124} + {{ 4 {bnn_N_Mux_2_2_3_1_3227_out1[1]}}, bnn_N_Mux_2_2_3_1_3227_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1859_out1 or bnn_Minus_2S_2S_1_3223_out1)
          begin :bnn_N_Mux_2_2_3_1_3241
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3241_out1 = bnn_Minus_2S_2S_1_3223_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3241_out1 = bnn_N_Mux_2_2_3_1_1859_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3243_in3 = {bnn_RightShift_64Sx8S_1S_1_3230_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3231_out1 or bnn_N_Mux_2_2_3_1_3243_in3)
          begin :bnn_N_Mux_2_2_3_1_3243
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3243_out1 = bnn_N_Mux_2_2_3_1_3231_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3243_out1 = bnn_N_Mux_2_2_3_1_3243_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3244_in1 = {s_reg_1041_stage1_slice[4:0], 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3244
         assign bnn_RightShift_64Sx8S_1S_1_3244_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3244_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3232_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3245
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3245_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3245_out1 = bnn_N_Mux_2_4_8_1_3232_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3246_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[44], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1974_out1 or bnn_N_Mux_2_2_3_1_1977_out1 or bnn_N_Mux_2_2_3_1_2089_out1 or bnn_N_Mux_2_4_8_1_3246_in3)
          begin :bnn_N_Mux_2_4_8_1_3246
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3246_out1 = bnn_N_Mux_2_2_3_1_1974_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3246_out1 = bnn_N_Mux_2_4_8_1_3246_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3246_out1 = bnn_N_Mux_2_2_3_1_1977_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3246_out1 = bnn_N_Mux_2_2_3_1_2089_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_41_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4446_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3247_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3247_in2 = {bnn_Mul_16Sx12S_19S_4_4446_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3247_in2 = {{ 5 {fixed_buffer_41_if_1_dout_wire[11]}}, fixed_buffer_41_if_1_dout_wire};
            end
         end

         // resource: mux_16bx3i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3234_out1[4:0] or gs_ctrl74)
          begin :drive_bnn_Add_17Sx16S_17S_1_3247_in1
            case (gs_ctrl74) 

               2'd1: begin
                  bnn_Add_17Sx16S_17S_1_3247_in1 = {{ 11 {s_reg_1138[4]}}, s_reg_1138[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_17Sx16S_17S_1_3247_in1 = s_reg_1138;
               end
               
               default: begin
                  bnn_Add_17Sx16S_17S_1_3247_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3234_out1[4]}}, bnn_Add_6Ux6U_6U_1_3234_out1[4:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3247
         assign bnn_Add_17Sx16S_17S_1_3247_out1 = bnn_Add_17Sx16S_17S_1_3247_in2 + {bnn_Add_17Sx16S_17S_1_3247_in1[15], bnn_Add_17Sx16S_17S_1_3247_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3236_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5014_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3248_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3248_in2 = bnn_Mod_6Ux32U_7U_4_5014_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3248_in2 = {bnn_Add_5Sx4S_6S_1_3236_out1[4], bnn_Add_5Sx4S_6S_1_3236_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1100[6:1] or bnn_N_Mux_2_2_3_4_3235_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3248_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3248_in1 = s_reg_1100[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3248_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3235_out1[1]}}, bnn_N_Mux_2_2_3_4_3235_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3248
         assign bnn_Add_6Ux6U_6U_1_3248_out1 = bnn_Add_6Ux6U_6U_1_3248_in2 + bnn_Add_6Ux6U_6U_1_3248_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1870_out1 or bnn_Minus_2S_2S_1_3237_out1)
          begin :bnn_N_Mux_2_2_3_4_3249
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3249_out1 = bnn_Minus_2S_2S_1_3237_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3249_out1 = bnn_N_Mux_2_2_3_1_1870_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3250
         assign bnn_Add_5Sx4S_6S_1_3250_out1 = {bnn_Add_5Sx4S_6S_1_3239_out1[4], bnn_Add_5Sx4S_6S_1_3239_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3238_out1[1]}}, bnn_N_Mux_2_2_3_1_3238_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3251
         assign bnn_Minus_2S_2S_1_3251_out1 = -bnn_N_Mux_2_2_3_1_1881_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1870_out1 or bnn_Minus_2S_2S_1_3237_out1)
          begin :bnn_N_Mux_2_2_3_1_3252
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3252_out1 = bnn_Minus_2S_2S_1_3237_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3252_out1 = bnn_N_Mux_2_2_3_1_1870_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3253
         assign bnn_Add_5Sx4S_6S_1_3253_out1 = {s_reg_1125[4], s_reg_1125} + {{ 4 {bnn_N_Mux_2_2_3_1_3241_out1[1]}}, bnn_N_Mux_2_2_3_1_3241_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1870_out1 or bnn_Minus_2S_2S_1_3237_out1)
          begin :bnn_N_Mux_2_2_3_1_3255
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3255_out1 = bnn_Minus_2S_2S_1_3237_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3255_out1 = bnn_N_Mux_2_2_3_1_1870_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3257
         assign bnn_Minus_2S_2S_1_3257_out1 = -bnn_N_Mux_2_2_3_1_1892_out1;

         assign bnn_N_Mux_2_2_3_1_3258_in3 = {bnn_RightShift_64Sx8S_1S_1_3244_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3245_out1 or bnn_N_Mux_2_2_3_1_3258_in3)
          begin :bnn_N_Mux_2_2_3_1_3258
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3258_out1 = bnn_N_Mux_2_2_3_1_3245_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3258_out1 = bnn_N_Mux_2_2_3_1_3258_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3259_in1 = {s_reg_1041_stage1_slice[4:0], 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3259
         assign bnn_RightShift_64Sx8S_1S_1_3259_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3259_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3246_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3260
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3260_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3260_out1 = bnn_N_Mux_2_4_8_1_3246_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3261_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[45], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1985_out1 or bnn_N_Mux_2_2_3_1_1988_out1 or bnn_N_Mux_2_2_3_1_2106_out1 or bnn_N_Mux_2_4_8_1_3261_in3)
          begin :bnn_N_Mux_2_4_8_1_3261
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3261_out1 = bnn_N_Mux_2_2_3_1_1985_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3261_out1 = bnn_N_Mux_2_4_8_1_3261_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3261_out1 = bnn_N_Mux_2_2_3_1_1988_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3261_out1 = bnn_N_Mux_2_2_3_1_2106_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_42_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4453_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3262_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3262_in2 = {bnn_Mul_16Sx12S_19S_4_4453_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3262_in2 = {{ 5 {fixed_buffer_42_if_1_dout_wire[11]}}, fixed_buffer_42_if_1_dout_wire};
            end
         end

         // resource: mux_16bx3i
         always @(s_reg_1138 or s_reg_1139 or bnn_Add_6Ux6U_6U_1_3248_out1[4:0] or gs_ctrl74)
          begin :drive_bnn_Add_17Sx16S_17S_1_3262_in1
            case (gs_ctrl74) 

               2'd1: begin
                  bnn_Add_17Sx16S_17S_1_3262_in1 = {{ 11 {s_reg_1139[4]}}, s_reg_1139};
               end
               
               2'd2: begin
                  bnn_Add_17Sx16S_17S_1_3262_in1 = s_reg_1138;
               end
               
               default: begin
                  bnn_Add_17Sx16S_17S_1_3262_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3248_out1[4]}}, bnn_Add_6Ux6U_6U_1_3248_out1[4:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3262
         assign bnn_Add_17Sx16S_17S_1_3262_out1 = bnn_Add_17Sx16S_17S_1_3262_in2 + {bnn_Add_17Sx16S_17S_1_3262_in1[15], bnn_Add_17Sx16S_17S_1_3262_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3250_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5015_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3263_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3263_in2 = bnn_Mod_6Ux32U_7U_4_5015_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3263_in2 = {bnn_Add_5Sx4S_6S_1_3250_out1[4], bnn_Add_5Sx4S_6S_1_3250_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1090[6:1] or bnn_N_Mux_2_2_3_4_3249_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3263_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3263_in1 = s_reg_1090[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3263_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3249_out1[1]}}, bnn_N_Mux_2_2_3_4_3249_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3263
         assign bnn_Add_6Ux6U_6U_1_3263_out1 = bnn_Add_6Ux6U_6U_1_3263_in2 + bnn_Add_6Ux6U_6U_1_3263_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1881_out1 or bnn_Minus_2S_2S_1_3251_out1)
          begin :bnn_N_Mux_2_2_3_1_3264
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3264_out1 = bnn_Minus_2S_2S_1_3251_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3264_out1 = bnn_N_Mux_2_2_3_1_1881_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3265
         assign bnn_Add_5Sx4S_6S_1_3265_out1 = {bnn_Add_5Sx4S_6S_1_3253_out1[4], bnn_Add_5Sx4S_6S_1_3253_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3252_out1[1]}}, bnn_N_Mux_2_2_3_1_3252_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1881_out1 or bnn_Minus_2S_2S_1_3251_out1)
          begin :bnn_N_Mux_2_2_3_1_3267
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3267_out1 = bnn_Minus_2S_2S_1_3251_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3267_out1 = bnn_N_Mux_2_2_3_1_1881_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3268
         assign bnn_Add_5Sx4S_6S_1_3268_out1 = {s_reg_1126[4], s_reg_1126} + {{ 4 {bnn_N_Mux_2_2_3_1_3255_out1[1]}}, bnn_N_Mux_2_2_3_1_3255_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1881_out1 or bnn_Minus_2S_2S_1_3251_out1)
          begin :bnn_N_Mux_2_2_3_4_3270
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3270_out1 = bnn_Minus_2S_2S_1_3251_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3270_out1 = bnn_N_Mux_2_2_3_1_1881_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3271
         assign bnn_Minus_2S_2S_4_3271_out1 = -bnn_N_Mux_2_2_3_1_1903_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1892_out1 or bnn_Minus_2S_2S_1_3257_out1)
          begin :bnn_N_Mux_2_2_3_4_3272
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3272_out1 = bnn_Minus_2S_2S_1_3257_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3272_out1 = bnn_N_Mux_2_2_3_1_1892_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3273
         assign bnn_Minus_2S_2S_1_3273_out1 = -bnn_N_Mux_2_2_3_1_2167_out1;

         assign bnn_N_Mux_2_2_3_1_3274_in3 = {bnn_RightShift_64Sx8S_1S_1_3259_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3260_out1 or bnn_N_Mux_2_2_3_1_3274_in3)
          begin :bnn_N_Mux_2_2_3_1_3274
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3274_out1 = bnn_N_Mux_2_2_3_1_3260_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3274_out1 = bnn_N_Mux_2_2_3_1_3274_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3275_in1 = {s_reg_1041_stage1_slice[4:0], 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3275
         assign bnn_RightShift_64Sx8S_1S_1_3275_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3275_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3261_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3276
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3276_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3276_out1 = bnn_N_Mux_2_4_8_1_3261_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3277_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[46], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_1996_out1 or bnn_N_Mux_2_2_3_1_1999_out1 or bnn_N_Mux_2_2_3_1_2123_out1 or bnn_N_Mux_2_4_8_1_3277_in3)
          begin :bnn_N_Mux_2_4_8_1_3277
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3277_out1 = bnn_N_Mux_2_2_3_1_1996_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3277_out1 = bnn_N_Mux_2_4_8_1_3277_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3277_out1 = bnn_N_Mux_2_2_3_1_1999_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3277_out1 = bnn_N_Mux_2_2_3_1_2123_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_43_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4440_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3278_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3278_in2 = {bnn_Mul_16Sx12S_19S_4_4440_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3278_in2 = {{ 5 {fixed_buffer_43_if_1_dout_wire[11]}}, fixed_buffer_43_if_1_dout_wire};
            end
         end

         // resource: mux_16bx3i
         always @(s_reg_1138 or s_reg_1140 or bnn_Add_6Ux6U_6U_1_3263_out1[4:0] or gs_ctrl74)
          begin :drive_bnn_Add_17Sx16S_17S_1_3278_in1
            case (gs_ctrl74) 

               2'd1: begin
                  bnn_Add_17Sx16S_17S_1_3278_in1 = {{ 11 {s_reg_1140[4]}}, s_reg_1140};
               end
               
               2'd2: begin
                  bnn_Add_17Sx16S_17S_1_3278_in1 = s_reg_1138;
               end
               
               default: begin
                  bnn_Add_17Sx16S_17S_1_3278_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3263_out1[4]}}, bnn_Add_6Ux6U_6U_1_3263_out1[4:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3278
         assign bnn_Add_17Sx16S_17S_1_3278_out1 = bnn_Add_17Sx16S_17S_1_3278_in2 + {bnn_Add_17Sx16S_17S_1_3278_in1[15], bnn_Add_17Sx16S_17S_1_3278_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3265_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5016_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3279_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3279_in2 = bnn_Mod_6Ux32U_7U_4_5016_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3279_in2 = {bnn_Add_5Sx4S_6S_1_3265_out1[4], bnn_Add_5Sx4S_6S_1_3265_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1092[6:1] or bnn_N_Mux_2_2_3_1_3264_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3279_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3279_in1 = s_reg_1092[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3279_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3264_out1[1]}}, bnn_N_Mux_2_2_3_1_3264_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3279
         assign bnn_Add_6Ux6U_6U_1_3279_out1 = bnn_Add_6Ux6U_6U_1_3279_in2 + bnn_Add_6Ux6U_6U_1_3279_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1892_out1 or bnn_Minus_2S_2S_1_3257_out1)
          begin :bnn_N_Mux_2_2_3_1_3280
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3280_out1 = bnn_Minus_2S_2S_1_3257_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3280_out1 = bnn_N_Mux_2_2_3_1_1892_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3281
         assign bnn_Add_5Sx4S_6S_1_3281_out1 = {bnn_Add_5Sx4S_6S_1_3268_out1[4], bnn_Add_5Sx4S_6S_1_3268_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3267_out1[1]}}, bnn_N_Mux_2_2_3_1_3267_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1892_out1 or bnn_Minus_2S_2S_1_3257_out1)
          begin :bnn_N_Mux_2_2_3_4_3283
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3283_out1 = bnn_Minus_2S_2S_1_3257_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3283_out1 = bnn_N_Mux_2_2_3_1_1892_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3284
         assign bnn_Add_5Sx4S_6S_1_3284_out1 = {s_reg_1127[4], s_reg_1127} + {{ 4 {bnn_N_Mux_2_2_3_4_3270_out1[1]}}, bnn_N_Mux_2_2_3_4_3270_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3285
         assign bnn_Minus_2S_2S_4_3285_out1 = -bnn_N_Mux_2_2_3_1_2155_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1903_out1 or bnn_Minus_2S_2S_4_3271_out1)
          begin :bnn_N_Mux_2_2_3_4_3286
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3286_out1 = bnn_Minus_2S_2S_4_3271_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3286_out1 = bnn_N_Mux_2_2_3_1_1903_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3287
         assign bnn_Add_5Sx4S_6S_1_3287_out1 = {s_reg_1128[4], s_reg_1128} + {{ 4 {bnn_N_Mux_2_2_3_4_3272_out1[1]}}, bnn_N_Mux_2_2_3_4_3272_out1};

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3288
         assign bnn_Minus_2S_2S_4_3288_out1 = -bnn_N_Mux_2_2_3_1_1924_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2167_out1 or bnn_Minus_2S_2S_1_3273_out1)
          begin :bnn_N_Mux_2_2_3_4_3289
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3289_out1 = bnn_Minus_2S_2S_1_3273_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3289_out1 = bnn_N_Mux_2_2_3_1_2167_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3290_in3 = {bnn_RightShift_64Sx8S_1S_1_3275_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3276_out1 or bnn_N_Mux_2_2_3_1_3290_in3)
          begin :bnn_N_Mux_2_2_3_1_3290
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3290_out1 = bnn_N_Mux_2_2_3_1_3276_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3290_out1 = bnn_N_Mux_2_2_3_1_3290_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3291_in1 = {s_reg_1041_stage1_slice[4:0], 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3291
         assign bnn_RightShift_64Sx8S_1S_1_3291_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3291_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3277_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3292
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3292_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3292_out1 = bnn_N_Mux_2_4_8_1_3277_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3293_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[47], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2007_out1 or bnn_N_Mux_2_2_3_1_2010_out1 or bnn_N_Mux_2_2_3_1_2140_out1 or bnn_N_Mux_2_4_8_1_3293_in3)
          begin :bnn_N_Mux_2_4_8_1_3293
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3293_out1 = bnn_N_Mux_2_2_3_1_2007_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3293_out1 = bnn_N_Mux_2_4_8_1_3293_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3293_out1 = bnn_N_Mux_2_2_3_1_2010_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3293_out1 = bnn_N_Mux_2_2_3_1_2140_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2205_out1 or bnn_N_Mux_2_2_3_1_2208_out1 or bnn_N_Mux_2_2_3_1_2214_out1 or bnn_N_Mux_3_2_6_4_1640_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3294
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3294_out1 = bnn_N_Mux_2_2_3_1_2205_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3294_out1 = bnn_N_Mux_3_2_6_4_1640_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3294_out1 = bnn_N_Mux_2_2_3_1_2208_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3294_out1 = bnn_N_Mux_2_2_3_1_2214_out1;
               end
               
            endcase

         end

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3295
         assign bnn_RightShift_64Sx8S_1S_4_3295_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_Sub_8Sx2S_8S_4_1610_out1[5:0];

         // resource: mux_17bx2i
         always @(fixed_buffer_44_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4462_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3296_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3296_in2 = {bnn_Mul_16Sx12S_19S_4_4462_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3296_in2 = {{ 5 {fixed_buffer_44_if_1_dout_wire[11]}}, fixed_buffer_44_if_1_dout_wire};
            end
         end

         // resource: mux_16bx3i
         always @(s_reg_1138 or s_reg_1141 or bnn_Add_6Ux6U_6U_1_3279_out1[4:0] or gs_ctrl74)
          begin :drive_bnn_Add_17Sx16S_17S_1_3296_in1
            case (gs_ctrl74) 

               2'd1: begin
                  bnn_Add_17Sx16S_17S_1_3296_in1 = {{ 11 {s_reg_1141[4]}}, s_reg_1141};
               end
               
               2'd2: begin
                  bnn_Add_17Sx16S_17S_1_3296_in1 = s_reg_1138;
               end
               
               default: begin
                  bnn_Add_17Sx16S_17S_1_3296_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3279_out1[4]}}, bnn_Add_6Ux6U_6U_1_3279_out1[4:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3296
         assign bnn_Add_17Sx16S_17S_1_3296_out1 = bnn_Add_17Sx16S_17S_1_3296_in2 + {bnn_Add_17Sx16S_17S_1_3296_in1[15], bnn_Add_17Sx16S_17S_1_3296_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3281_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5017_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3297_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3297_in2 = bnn_Mod_6Ux32U_7U_4_5017_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3297_in2 = {bnn_Add_5Sx4S_6S_1_3281_out1[4], bnn_Add_5Sx4S_6S_1_3281_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1089[6:1] or bnn_N_Mux_2_2_3_1_3280_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3297_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3297_in1 = s_reg_1089[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3297_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3280_out1[1]}}, bnn_N_Mux_2_2_3_1_3280_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3297
         assign bnn_Add_6Ux6U_6U_1_3297_out1 = bnn_Add_6Ux6U_6U_1_3297_in2 + bnn_Add_6Ux6U_6U_1_3297_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1903_out1 or bnn_Minus_2S_2S_4_3271_out1)
          begin :bnn_N_Mux_2_2_3_4_3298
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3298_out1 = bnn_Minus_2S_2S_4_3271_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3298_out1 = bnn_N_Mux_2_2_3_1_1903_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3299
         assign bnn_Add_5Sx4S_6S_1_3299_out1 = {bnn_Add_5Sx4S_6S_1_3284_out1[4], bnn_Add_5Sx4S_6S_1_3284_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3283_out1[1]}}, bnn_N_Mux_2_2_3_4_3283_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2155_out1 or bnn_Minus_2S_2S_4_3285_out1)
          begin :bnn_N_Mux_2_2_3_4_3301
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3301_out1 = bnn_Minus_2S_2S_4_3285_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3301_out1 = bnn_N_Mux_2_2_3_1_2155_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3302
         assign bnn_Add_5Sx4S_6S_1_3302_out1 = {bnn_Add_5Sx4S_6S_1_3287_out1[4], bnn_Add_5Sx4S_6S_1_3287_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3286_out1[1]}}, bnn_N_Mux_2_2_3_4_3286_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3303
         assign bnn_Minus_2S_2S_1_3303_out1 = -bnn_N_Mux_2_2_3_1_1935_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1924_out1 or bnn_Minus_2S_2S_4_3288_out1)
          begin :bnn_N_Mux_2_2_3_4_3304
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3304_out1 = bnn_Minus_2S_2S_4_3288_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3304_out1 = bnn_N_Mux_2_2_3_1_1924_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3305
         assign bnn_Add_5Sx4S_6S_1_3305_out1 = {s_reg_1129[4], s_reg_1129} + {{ 4 {bnn_N_Mux_2_2_3_4_3289_out1[1]}}, bnn_N_Mux_2_2_3_4_3289_out1};

         assign bnn_N_Mux_2_2_3_1_3306_in3 = {bnn_RightShift_64Sx8S_1S_1_3291_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3292_out1 or bnn_N_Mux_2_2_3_1_3306_in3)
          begin :bnn_N_Mux_2_2_3_1_3306
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3306_out1 = bnn_N_Mux_2_2_3_1_3292_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3306_out1 = bnn_N_Mux_2_2_3_1_3306_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3307_in1 = {s_reg_1041_stage1_slice[4:0], 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3307
         assign bnn_RightShift_64Sx8S_1S_1_3307_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3307_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3293_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3308
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3308_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3308_out1 = bnn_N_Mux_2_4_8_1_3293_out1;
            end
         end

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2187_out1 or bnn_N_Mux_2_2_3_1_2190_out1 or bnn_N_Mux_2_2_3_1_2196_out1 or bnn_N_Mux_3_2_6_1_1639_out1_slice)
          begin :bnn_N_Mux_2_4_8_1_3309
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3309_out1 = bnn_N_Mux_2_2_3_1_2187_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3309_out1 = bnn_N_Mux_3_2_6_1_1639_out1_slice;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3309_out1 = bnn_N_Mux_2_2_3_1_2190_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3309_out1 = bnn_N_Mux_2_2_3_1_2196_out1;
               end
               
            endcase

         end

         assign bnn_RightShift_64Sx8S_1S_1_3310_in1 = {s_reg_1109, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3310
         assign bnn_RightShift_64Sx8S_1S_1_3310_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3310_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3294_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3311
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3311_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3311_out1 = bnn_N_Mux_2_4_8_4_3294_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_4_3312_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_4_3295_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(bnn_N_Mux_3_2_6_4_3312_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_4_3312
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_4_3312_out1_slice = bnn_N_Mux_3_2_6_4_3312_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_3312_out1_slice = 2'd0;
            end
         end

         assign bnn_N_Mux_2_4_8_1_3313_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[48], 1'b1};

         // resource: bnn_N_Mux_2_4_8_1
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2018_out1 or bnn_N_Mux_2_2_3_1_2021_out1 or bnn_N_Mux_2_2_3_1_2027_out1 or bnn_N_Mux_2_4_8_1_3313_in3)
          begin :bnn_N_Mux_2_4_8_1_3313
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_1_3313_out1 = bnn_N_Mux_2_2_3_1_2018_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_1_3313_out1 = bnn_N_Mux_2_4_8_1_3313_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_1_3313_out1 = bnn_N_Mux_2_2_3_1_2021_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_1_3313_out1 = bnn_N_Mux_2_2_3_1_2027_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_45_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4436_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3314_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3314_in2 = {bnn_Mul_16Sx12S_19S_4_4436_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3314_in2 = {{ 5 {fixed_buffer_45_if_1_dout_wire[11]}}, fixed_buffer_45_if_1_dout_wire};
            end
         end

         // resource: mux_16bx3i
         always @(s_reg_1138 or s_reg_1142 or bnn_Add_6Ux6U_6U_1_3297_out1[4:0] or gs_ctrl74)
          begin :drive_bnn_Add_17Sx16S_17S_1_3314_in1
            case (gs_ctrl74) 

               2'd1: begin
                  bnn_Add_17Sx16S_17S_1_3314_in1 = {{ 11 {s_reg_1142[4]}}, s_reg_1142};
               end
               
               2'd2: begin
                  bnn_Add_17Sx16S_17S_1_3314_in1 = s_reg_1138;
               end
               
               default: begin
                  bnn_Add_17Sx16S_17S_1_3314_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3297_out1[4]}}, bnn_Add_6Ux6U_6U_1_3297_out1[4:0]};
               end
               
            endcase

         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3314
         assign bnn_Add_17Sx16S_17S_1_3314_out1 = bnn_Add_17Sx16S_17S_1_3314_in2 + {bnn_Add_17Sx16S_17S_1_3314_in1[15], bnn_Add_17Sx16S_17S_1_3314_in1};

         // resource: mux_6bx3i
         always @(s_reg_1047 or bnn_Add_5Sx4S_6S_1_3299_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4998_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3315_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3315_in2 = {s_reg_1047[4], s_reg_1047};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3315_in2 = bnn_Mod_6Ux32U_7U_4_4998_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3315_in2 = {bnn_Add_5Sx4S_6S_1_3299_out1[4], bnn_Add_5Sx4S_6S_1_3299_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1025[6:1] or s_reg_1115[1:0] or bnn_N_Mux_2_2_3_4_3298_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3315_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3315_in1 = {{ 4 {s_reg_1115[1]}}, s_reg_1115[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3315_in1 = s_reg_1025[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3315_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3298_out1[1]}}, bnn_N_Mux_2_2_3_4_3298_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3315
         assign bnn_Add_6Ux6U_6U_1_3315_out1 = bnn_Add_6Ux6U_6U_1_3315_in2 + bnn_Add_6Ux6U_6U_1_3315_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1924_out1 or bnn_Minus_2S_2S_4_3288_out1)
          begin :bnn_N_Mux_2_2_3_4_3317
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3317_out1 = bnn_Minus_2S_2S_4_3288_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3317_out1 = bnn_N_Mux_2_2_3_1_1924_out1;
            end
         end

         // resource: mux_6bx3i
         always @(s_reg_871 or bnn_Add_5Sx4S_6S_1_3302_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4999_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3319_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3319_in2 = {s_reg_871[4], s_reg_871};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3319_in2 = bnn_Mod_6Ux32U_7U_4_4999_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3319_in2 = {bnn_Add_5Sx4S_6S_1_3302_out1[4], bnn_Add_5Sx4S_6S_1_3302_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1091[6:1] or s_reg_1116[1:0] or bnn_N_Mux_2_2_3_4_3301_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3319_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3319_in1 = {{ 4 {s_reg_1116[1]}}, s_reg_1116[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3319_in1 = s_reg_1091[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3319_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3301_out1[1]}}, bnn_N_Mux_2_2_3_4_3301_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3319
         assign bnn_Add_6Ux6U_6U_1_3319_out1 = bnn_Add_6Ux6U_6U_1_3319_in2 + bnn_Add_6Ux6U_6U_1_3319_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1935_out1 or bnn_Minus_2S_2S_1_3303_out1)
          begin :bnn_N_Mux_2_2_3_4_3320
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3320_out1 = bnn_Minus_2S_2S_1_3303_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3320_out1 = bnn_N_Mux_2_2_3_1_1935_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3321
         assign bnn_Add_5Sx4S_6S_1_3321_out1 = {bnn_Add_5Sx4S_6S_1_3305_out1[4], bnn_Add_5Sx4S_6S_1_3305_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3304_out1[1]}}, bnn_N_Mux_2_2_3_4_3304_out1};

         assign bnn_N_Mux_2_2_3_1_3322_in3 = {bnn_RightShift_64Sx8S_1S_1_3307_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3308_out1 or bnn_N_Mux_2_2_3_1_3322_in3)
          begin :bnn_N_Mux_2_2_3_1_3322
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3322_out1 = bnn_N_Mux_2_2_3_1_3308_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3322_out1 = bnn_N_Mux_2_2_3_1_3322_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3309_out1 or s_reg_1057_stage1)
          begin :bnn_N_Mux_2_2_3_1_3323
            if (s_reg_1057_stage1) begin
               bnn_N_Mux_2_2_3_1_3323_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3323_out1 = bnn_N_Mux_2_4_8_1_3309_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_1_3324_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_1_3310_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_1
         always @(bnn_N_Mux_3_2_6_1_3324_in2[1:0] or s_reg_1088_stage1)
          begin :bnn_N_Mux_3_2_6_1_3324
            if (s_reg_1088_stage1) begin
               bnn_N_Mux_3_2_6_1_3324_out1_slice = bnn_N_Mux_3_2_6_1_3324_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_1_3324_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3311_out1 or bnn_N_Mux_3_2_6_4_3312_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_3325
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3325_out1 = bnn_N_Mux_2_2_3_4_3311_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3325_out1 = bnn_N_Mux_3_2_6_4_3312_out1_slice;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_1_3326_in1 = {s_reg_1058_stage1_slice[4:0], 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_1  instance: bnn_RightShift_64Sx8S_1S_1_3326
         assign bnn_RightShift_64Sx8S_1S_1_3326_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_1_3326_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_N_Mux_2_4_8_1_3313_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_1_3327
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_1_3327_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3327_out1 = bnn_N_Mux_2_4_8_1_3313_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3328_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[49], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2035_out1 or bnn_N_Mux_2_2_3_1_2038_out1 or bnn_N_Mux_2_2_3_1_2044_out1 or bnn_N_Mux_2_4_8_4_3328_in3)
          begin :bnn_N_Mux_2_4_8_4_3328
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3328_out1 = bnn_N_Mux_2_2_3_1_2035_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3328_out1 = bnn_N_Mux_2_4_8_4_3328_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3328_out1 = bnn_N_Mux_2_2_3_1_2038_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3328_out1 = bnn_N_Mux_2_2_3_1_2044_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_46_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4551_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3329_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3329_in2 = {bnn_Mul_16Sx12S_19S_4_4551_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3329_in2 = {{ 5 {fixed_buffer_46_if_1_dout_wire[11]}}, fixed_buffer_46_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3315_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3329_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3329_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3329_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3315_out1[4]}}, bnn_Add_6Ux6U_6U_1_3315_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3329
         assign bnn_Add_17Sx16S_17S_1_3329_out1 = bnn_Add_17Sx16S_17S_1_3329_in2 + {bnn_Add_17Sx16S_17S_1_3329_in1[15], bnn_Add_17Sx16S_17S_1_3329_in1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3330
         assign bnn_Minus_2S_2S_1_3330_out1 = -bnn_N_Mux_2_2_3_1_1946_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1935_out1 or bnn_Minus_2S_2S_1_3303_out1)
          begin :bnn_N_Mux_2_2_3_4_3331
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3331_out1 = bnn_Minus_2S_2S_1_3303_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3331_out1 = bnn_N_Mux_2_2_3_1_1935_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3332
         assign bnn_Add_5Sx4S_6S_1_3332_out1 = {s_reg_1131[4], s_reg_1131} + {{ 4 {bnn_N_Mux_2_2_3_4_3317_out1[1]}}, bnn_N_Mux_2_2_3_4_3317_out1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1935_out1 or bnn_Minus_2S_2S_1_3303_out1)
          begin :bnn_N_Mux_2_2_3_4_3334
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3334_out1 = bnn_Minus_2S_2S_1_3303_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3334_out1 = bnn_N_Mux_2_2_3_1_1935_out1;
            end
         end

         // resource: mux_6bx3i
         always @(s_reg_1091[4:0] or bnn_Add_5Sx4S_6S_1_3321_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4989_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3336_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3336_in2 = {s_reg_1091[4], s_reg_1091[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3336_in2 = bnn_Mod_6Ux32U_7U_4_4989_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3336_in2 = {bnn_Add_5Sx4S_6S_1_3321_out1[4], bnn_Add_5Sx4S_6S_1_3321_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1106[6:1] or s_reg_1117[1:0] or bnn_N_Mux_2_2_3_4_3320_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3336_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3336_in1 = {{ 4 {s_reg_1117[1]}}, s_reg_1117[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3336_in1 = s_reg_1106[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3336_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3320_out1[1]}}, bnn_N_Mux_2_2_3_4_3320_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3336
         assign bnn_Add_6Ux6U_6U_1_3336_out1 = bnn_Add_6Ux6U_6U_1_3336_in2 + bnn_Add_6Ux6U_6U_1_3336_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1581_out1 or bnn_N_Mux_2_2_3_1_3323_out1 or bnn_N_Mux_3_2_6_1_3324_out1_slice)
          begin :bnn_N_Mux_2_2_3_1_3337
            if (bnn_Or_1Sx1U_1S_4_1581_out1) begin
               bnn_N_Mux_2_2_3_1_3337_out1 = bnn_N_Mux_2_2_3_1_3323_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3337_out1 = bnn_N_Mux_3_2_6_1_3324_out1_slice;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3338_in3 = {bnn_RightShift_64Sx8S_1S_1_3326_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_1_3327_out1 or bnn_N_Mux_2_2_3_1_3338_in3)
          begin :bnn_N_Mux_2_2_3_1_3338
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_1_3338_out1 = bnn_N_Mux_2_2_3_1_3327_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3338_out1 = bnn_N_Mux_2_2_3_1_3338_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3339_in1 = {s_reg_1058_stage1_slice[4:0], 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3339
         assign bnn_RightShift_64Sx8S_1S_4_3339_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3339_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3328_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3340
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3340_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3340_out1 = bnn_N_Mux_2_4_8_4_3328_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3341_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[50], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2052_out1 or bnn_N_Mux_2_2_3_1_2055_out1 or bnn_N_Mux_2_2_3_1_2061_out1 or bnn_N_Mux_2_4_8_4_3341_in3)
          begin :bnn_N_Mux_2_4_8_4_3341
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3341_out1 = bnn_N_Mux_2_2_3_1_2052_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3341_out1 = bnn_N_Mux_2_4_8_4_3341_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3341_out1 = bnn_N_Mux_2_2_3_1_2055_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3341_out1 = bnn_N_Mux_2_2_3_1_2061_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_47_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4561_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3342_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3342_in2 = {bnn_Mul_16Sx12S_19S_4_4561_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3342_in2 = {{ 5 {fixed_buffer_47_if_1_dout_wire[11]}}, fixed_buffer_47_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3319_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3342_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3342_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3342_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3319_out1[4]}}, bnn_Add_6Ux6U_6U_1_3319_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3342
         assign bnn_Add_17Sx16S_17S_1_3342_out1 = bnn_Add_17Sx16S_17S_1_3342_in2 + {bnn_Add_17Sx16S_17S_1_3342_in1[15], bnn_Add_17Sx16S_17S_1_3342_in1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_1946_out1 or bnn_Minus_2S_2S_1_3330_out1)
          begin :bnn_N_Mux_2_2_3_4_3343
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3343_out1 = bnn_Minus_2S_2S_1_3330_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3343_out1 = bnn_N_Mux_2_2_3_1_1946_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3344
         assign bnn_Add_5Sx4S_6S_1_3344_out1 = {bnn_Add_5Sx4S_6S_1_3332_out1[4], bnn_Add_5Sx4S_6S_1_3332_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3331_out1[1]}}, bnn_N_Mux_2_2_3_4_3331_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3345
         assign bnn_Minus_2S_2S_1_3345_out1 = -bnn_N_Mux_2_2_3_1_1957_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_1946_out1 or bnn_Minus_2S_2S_1_3330_out1)
          begin :bnn_N_Mux_2_2_3_4_3346
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3346_out1 = bnn_Minus_2S_2S_1_3330_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3346_out1 = bnn_N_Mux_2_2_3_1_1946_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3347
         assign bnn_Add_5Sx4S_6S_1_3347_out1 = {s_reg_1132[4], s_reg_1132} + {{ 4 {bnn_N_Mux_2_2_3_4_3334_out1[1]}}, bnn_N_Mux_2_2_3_4_3334_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1946_out1 or bnn_Minus_2S_2S_1_3330_out1)
          begin :bnn_N_Mux_2_2_3_1_3349
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3349_out1 = bnn_Minus_2S_2S_1_3330_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3349_out1 = bnn_N_Mux_2_2_3_1_1946_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3351_in3 = {bnn_RightShift_64Sx8S_1S_4_3339_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3340_out1 or bnn_N_Mux_2_2_3_4_3351_in3)
          begin :bnn_N_Mux_2_2_3_4_3351
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3351_out1 = bnn_N_Mux_2_2_3_4_3340_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3351_out1 = bnn_N_Mux_2_2_3_4_3351_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3341_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3353
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3353_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3353_out1 = bnn_N_Mux_2_4_8_4_3341_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3354_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[51], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2069_out1 or bnn_N_Mux_2_2_3_1_2072_out1 or bnn_N_Mux_2_2_3_1_2078_out1 or bnn_N_Mux_2_4_8_4_3354_in3)
          begin :bnn_N_Mux_2_4_8_4_3354
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3354_out1 = bnn_N_Mux_2_2_3_1_2069_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3354_out1 = bnn_N_Mux_2_4_8_4_3354_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3354_out1 = bnn_N_Mux_2_2_3_1_2072_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3354_out1 = bnn_N_Mux_2_2_3_1_2078_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_48_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4571_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3355_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3355_in2 = {bnn_Mul_16Sx12S_19S_4_4571_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3355_in2 = {{ 5 {fixed_buffer_48_if_1_dout_wire[11]}}, fixed_buffer_48_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3336_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3355_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3355_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3355_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3336_out1[4]}}, bnn_Add_6Ux6U_6U_1_3336_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3355
         assign bnn_Add_17Sx16S_17S_1_3355_out1 = bnn_Add_17Sx16S_17S_1_3355_in2 + {bnn_Add_17Sx16S_17S_1_3355_in1[15], bnn_Add_17Sx16S_17S_1_3355_in1};

         // resource: mux_6bx3i
         always @(s_reg_1095[4:0] or bnn_Add_5Sx4S_6S_1_3344_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5000_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3356_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3356_in2 = {s_reg_1095[4], s_reg_1095[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3356_in2 = bnn_Mod_6Ux32U_7U_4_5000_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3356_in2 = {bnn_Add_5Sx4S_6S_1_3344_out1[4], bnn_Add_5Sx4S_6S_1_3344_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1076[6:1] or s_reg_1120[1:0] or bnn_N_Mux_2_2_3_4_3343_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3356_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3356_in1 = {{ 4 {s_reg_1120[1]}}, s_reg_1120[1:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3356_in1 = s_reg_1076[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3356_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3343_out1[1]}}, bnn_N_Mux_2_2_3_4_3343_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3356
         assign bnn_Add_6Ux6U_6U_1_3356_out1 = bnn_Add_6Ux6U_6U_1_3356_in2 + bnn_Add_6Ux6U_6U_1_3356_in1;

         // resource: mux_2bx2i
         always @(s_reg_962 or bnn_N_Mux_2_2_3_1_1957_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3357_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3357_in3 = s_reg_962;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3357_in3 = bnn_N_Mux_2_2_3_1_1957_out1;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_Minus_2S_2S_1_1295_out1 or bnn_Minus_2S_2S_1_3345_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3357_in2
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3357_in2 = bnn_Minus_2S_2S_1_1295_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3357_in2 = bnn_Minus_2S_2S_1_3345_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_3357_in3 or bnn_N_Mux_2_2_3_1_3357_in2)
          begin :bnn_N_Mux_2_2_3_1_3357
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3357_out1 = bnn_N_Mux_2_2_3_1_3357_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3357_out1 = bnn_N_Mux_2_2_3_1_3357_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1097[4:0] or bnn_Add_5Sx4S_6S_1_3347_out1[4:0] or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3358_in2
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3358_in2 = s_reg_1097[4:0];
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3358_in2 = bnn_Add_5Sx4S_6S_1_3347_out1[4:0];
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_1121[1:0] or bnn_N_Mux_2_2_3_4_3346_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3358_in1
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3358_in1_slice = s_reg_1121[1:0];
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3358_in1_slice = bnn_N_Mux_2_2_3_4_3346_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3358
         assign bnn_Add_5Sx4S_6S_1_3358_out1 = {bnn_Add_5Sx4S_6S_1_3358_in2[4], bnn_Add_5Sx4S_6S_1_3358_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_3358_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_3358_in1_slice};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3359
         assign bnn_Minus_2S_2S_1_3359_out1 = -bnn_N_Mux_2_2_3_1_1968_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_3357_in3 or bnn_N_Mux_2_2_3_1_3357_in2)
          begin :bnn_N_Mux_2_2_3_1_3360
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3360_out1 = bnn_N_Mux_2_2_3_1_3357_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3360_out1 = bnn_N_Mux_2_2_3_1_3357_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1957_out1 or bnn_Minus_2S_2S_1_3345_out1)
          begin :bnn_N_Mux_2_2_3_1_3363
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3363_out1 = bnn_Minus_2S_2S_1_3345_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3363_out1 = bnn_N_Mux_2_2_3_1_1957_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_1_3365_in3 = {bnn_RightShift_64Sx8S_1S_1_228_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3353_out1 or bnn_N_Mux_2_2_3_1_3365_in3)
          begin :bnn_N_Mux_2_2_3_1_3365
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_1_3365_out1 = bnn_N_Mux_2_2_3_4_3353_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3365_out1 = bnn_N_Mux_2_2_3_1_3365_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3366_in1 = {s_reg_1058_stage1_slice[4:0], 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3366
         assign bnn_RightShift_64Sx8S_1S_4_3366_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3366_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3354_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3367
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3367_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3367_out1 = bnn_N_Mux_2_4_8_4_3354_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3368_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[52], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2086_out1 or bnn_N_Mux_2_2_3_1_2089_out1 or bnn_N_Mux_2_2_3_1_2095_out1 or bnn_N_Mux_2_4_8_4_3368_in3)
          begin :bnn_N_Mux_2_4_8_4_3368
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3368_out1 = bnn_N_Mux_2_2_3_1_2086_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3368_out1 = bnn_N_Mux_2_4_8_4_3368_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3368_out1 = bnn_N_Mux_2_2_3_1_2089_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3368_out1 = bnn_N_Mux_2_2_3_1_2095_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_49_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4580_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3369_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3369_in2 = {bnn_Mul_16Sx12S_19S_4_4580_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3369_in2 = {{ 5 {fixed_buffer_49_if_1_dout_wire[11]}}, fixed_buffer_49_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3356_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3369_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3369_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3369_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3356_out1[4]}}, bnn_Add_6Ux6U_6U_1_3356_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3369
         assign bnn_Add_17Sx16S_17S_1_3369_out1 = bnn_Add_17Sx16S_17S_1_3369_in2 + {bnn_Add_17Sx16S_17S_1_3369_in1[15], bnn_Add_17Sx16S_17S_1_3369_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3358_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5001_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3370_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3370_in2 = bnn_Mod_6Ux32U_7U_4_5001_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3370_in2 = {bnn_Add_5Sx4S_6S_1_3358_out1[4], bnn_Add_5Sx4S_6S_1_3358_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1070[6:1] or bnn_N_Mux_2_2_3_1_3357_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3370_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3370_in1 = s_reg_1070[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3370_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3357_out1[1]}}, bnn_N_Mux_2_2_3_1_3357_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3370
         assign bnn_Add_6Ux6U_6U_1_3370_out1 = bnn_Add_6Ux6U_6U_1_3370_in2 + bnn_Add_6Ux6U_6U_1_3370_in1;

         // resource: mux_2bx2i
         always @(s_reg_965 or bnn_N_Mux_2_2_3_1_1968_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3371_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3371_in3 = s_reg_965;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3371_in3 = bnn_N_Mux_2_2_3_1_1968_out1;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_Minus_2S_2S_1_1386_out1 or bnn_Minus_2S_2S_1_3359_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3371_in2
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3371_in2 = bnn_Minus_2S_2S_1_1386_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3371_in2 = bnn_Minus_2S_2S_1_3359_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_3371_in3 or bnn_N_Mux_2_2_3_1_3371_in2)
          begin :bnn_N_Mux_2_2_3_1_3371
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3371_out1 = bnn_N_Mux_2_2_3_1_3371_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3371_out1 = bnn_N_Mux_2_2_3_1_3371_in3;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3372
         assign bnn_Add_5Sx4S_6S_1_3372_out1 = {bnn_Add_6Ux6U_6U_1_206_out1[4], bnn_Add_6Ux6U_6U_1_206_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3360_out1[1]}}, bnn_N_Mux_2_2_3_1_3360_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3373
         assign bnn_Minus_2S_2S_1_3373_out1 = -bnn_N_Mux_2_2_3_1_1979_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_3371_in3 or bnn_N_Mux_2_2_3_1_3371_in2)
          begin :bnn_N_Mux_2_2_3_1_3374
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3374_out1 = bnn_N_Mux_2_2_3_1_3371_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3374_out1 = bnn_N_Mux_2_2_3_1_3371_in3;
            end
         end

         // resource: mux_6bx3i
         always @(s_reg_1134 or bnn_Add_5Sx3S_5S_1_209_out1 or bnn_N_Mux_6_2_12_4_4443_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3375_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3375_in2 = {bnn_Add_5Sx3S_5S_1_209_out1[4], bnn_Add_5Sx3S_5S_1_209_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3375_in2 = bnn_N_Mux_6_2_12_4_4443_out1;
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3375_in2 = {s_reg_1134[4], s_reg_1134};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(bnn_N_Mux_2_2_3_1_1454_out1 or bnn_N_Mux_2_2_3_1_3363_out1 or bnn_LeftShift_9Ux3U_7U_4_4442_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3375_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3375_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1454_out1[1]}}, bnn_N_Mux_2_2_3_1_1454_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3375_in1 = bnn_LeftShift_9Ux3U_7U_4_4442_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3375_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3363_out1[1]}}, bnn_N_Mux_2_2_3_1_3363_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3375
         assign bnn_Add_6Ux6U_6U_1_3375_out1 = bnn_Add_6Ux6U_6U_1_3375_in2 + bnn_Add_6Ux6U_6U_1_3375_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1968_out1 or bnn_Minus_2S_2S_1_3359_out1)
          begin :bnn_N_Mux_2_2_3_1_3377
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3377_out1 = bnn_Minus_2S_2S_1_3359_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3377_out1 = bnn_N_Mux_2_2_3_1_1968_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3379
         assign bnn_Minus_2S_2S_1_3379_out1 = -bnn_N_Mux_2_2_3_1_1990_out1;

         assign bnn_N_Mux_2_2_3_4_3380_in3 = {bnn_RightShift_64Sx8S_1S_4_3366_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3367_out1 or bnn_N_Mux_2_2_3_4_3380_in3)
          begin :bnn_N_Mux_2_2_3_4_3380
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3380_out1 = bnn_N_Mux_2_2_3_4_3367_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3380_out1 = bnn_N_Mux_2_2_3_4_3380_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3381_in1 = {s_reg_1058_stage1_slice[4:0], 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3381
         assign bnn_RightShift_64Sx8S_1S_4_3381_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3381_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3368_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3382
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3382_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3382_out1 = bnn_N_Mux_2_4_8_4_3368_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3383_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[53], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2103_out1 or bnn_N_Mux_2_2_3_1_2106_out1 or bnn_N_Mux_2_2_3_1_2112_out1 or bnn_N_Mux_2_4_8_4_3383_in3)
          begin :bnn_N_Mux_2_4_8_4_3383
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3383_out1 = bnn_N_Mux_2_2_3_1_2103_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3383_out1 = bnn_N_Mux_2_4_8_4_3383_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3383_out1 = bnn_N_Mux_2_2_3_1_2106_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3383_out1 = bnn_N_Mux_2_2_3_1_2112_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_50_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4589_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3384_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3384_in2 = {bnn_Mul_16Sx12S_19S_4_4589_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3384_in2 = {{ 5 {fixed_buffer_50_if_1_dout_wire[11]}}, fixed_buffer_50_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3370_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3384_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3384_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3384_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3370_out1[4]}}, bnn_Add_6Ux6U_6U_1_3370_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3384
         assign bnn_Add_17Sx16S_17S_1_3384_out1 = bnn_Add_17Sx16S_17S_1_3384_in2 + {bnn_Add_17Sx16S_17S_1_3384_in1[15], bnn_Add_17Sx16S_17S_1_3384_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3372_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5002_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3385_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3385_in2 = bnn_Mod_6Ux32U_7U_4_5002_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3385_in2 = {bnn_Add_5Sx4S_6S_1_3372_out1[4], bnn_Add_5Sx4S_6S_1_3372_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1068[6:1] or bnn_N_Mux_2_2_3_1_3371_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3385_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3385_in1 = s_reg_1068[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3385_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3371_out1[1]}}, bnn_N_Mux_2_2_3_1_3371_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3385
         assign bnn_Add_6Ux6U_6U_1_3385_out1 = bnn_Add_6Ux6U_6U_1_3385_in2 + bnn_Add_6Ux6U_6U_1_3385_in1;

         // resource: mux_2bx2i
         always @(s_reg_968 or bnn_N_Mux_2_2_3_1_1979_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3386_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3386_in3 = s_reg_968;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3386_in3 = bnn_N_Mux_2_2_3_1_1979_out1;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_Minus_2S_2S_1_1397_out1 or bnn_Minus_2S_2S_1_3373_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3386_in2
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3386_in2 = bnn_Minus_2S_2S_1_1397_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3386_in2 = bnn_Minus_2S_2S_1_3373_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_3386_in3 or bnn_N_Mux_2_2_3_1_3386_in2)
          begin :bnn_N_Mux_2_2_3_1_3386
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3386_out1 = bnn_N_Mux_2_2_3_1_3386_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3386_out1 = bnn_N_Mux_2_2_3_1_3386_in3;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3387
         assign bnn_Add_5Sx4S_6S_1_3387_out1 = {bnn_Add_6Ux6U_6U_1_3375_out1[4], bnn_Add_6Ux6U_6U_1_3375_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3374_out1[1]}}, bnn_N_Mux_2_2_3_1_3374_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_3386_in3 or bnn_N_Mux_2_2_3_1_3386_in2)
          begin :bnn_N_Mux_2_2_3_1_3389
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3389_out1 = bnn_N_Mux_2_2_3_1_3386_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3389_out1 = bnn_N_Mux_2_2_3_1_3386_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1135 or bnn_Add_4Sx2S_5S_1_2289_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3390_in2
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3390_in2 = bnn_Add_4Sx2S_5S_1_2289_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3390_in2 = s_reg_1135;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_N_Mux_2_2_3_1_3377_out1 or bnn_N_Mux_2_2_3_1_3730_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3390_in1
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3390_in1_slice = bnn_N_Mux_2_2_3_1_3730_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3390_in1_slice = bnn_N_Mux_2_2_3_1_3377_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3390
         assign bnn_Add_5Sx4S_6S_1_3390_out1 = {bnn_Add_5Sx4S_6S_1_3390_in2[4], bnn_Add_5Sx4S_6S_1_3390_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_3390_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_3390_in1_slice};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1979_out1 or bnn_Minus_2S_2S_1_3373_out1)
          begin :bnn_N_Mux_2_2_3_1_3392
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3392_out1 = bnn_Minus_2S_2S_1_3373_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3392_out1 = bnn_N_Mux_2_2_3_1_1979_out1;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_974 or bnn_N_Mux_2_2_3_1_2001_out1 or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_4_3393_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_4_3393_in1 = s_reg_974;
            end
            else begin
               bnn_Minus_2S_2S_4_3393_in1 = bnn_N_Mux_2_2_3_1_2001_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3393
         assign bnn_Minus_2S_2S_4_3393_out1 = -bnn_Minus_2S_2S_4_3393_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_1990_out1 or bnn_Minus_2S_2S_1_3379_out1)
          begin :bnn_N_Mux_2_2_3_1_3394
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3394_out1 = bnn_Minus_2S_2S_1_3379_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3394_out1 = bnn_N_Mux_2_2_3_1_1990_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3395
         assign bnn_Minus_2S_2S_4_3395_out1 = -bnn_N_Mux_2_2_3_1_2199_out1;

         assign bnn_N_Mux_2_2_3_4_3396_in3 = {bnn_RightShift_64Sx8S_1S_4_3381_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3382_out1 or bnn_N_Mux_2_2_3_4_3396_in3)
          begin :bnn_N_Mux_2_2_3_4_3396
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3396_out1 = bnn_N_Mux_2_2_3_4_3382_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3396_out1 = bnn_N_Mux_2_2_3_4_3396_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3397_in1 = {s_reg_1058_stage1_slice[4:0], 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3397
         assign bnn_RightShift_64Sx8S_1S_4_3397_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3397_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3383_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3398
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3398_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3398_out1 = bnn_N_Mux_2_4_8_4_3383_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3399_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[54], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2120_out1 or bnn_N_Mux_2_2_3_1_2123_out1 or bnn_N_Mux_2_2_3_1_2129_out1 or bnn_N_Mux_2_4_8_4_3399_in3)
          begin :bnn_N_Mux_2_4_8_4_3399
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3399_out1 = bnn_N_Mux_2_2_3_1_2120_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3399_out1 = bnn_N_Mux_2_4_8_4_3399_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3399_out1 = bnn_N_Mux_2_2_3_1_2123_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3399_out1 = bnn_N_Mux_2_2_3_1_2129_out1;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_51_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4598_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3400_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3400_in2 = {bnn_Mul_16Sx12S_19S_4_4598_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3400_in2 = {{ 5 {fixed_buffer_51_if_1_dout_wire[11]}}, fixed_buffer_51_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3385_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3400_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3400_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3400_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3385_out1[4]}}, bnn_Add_6Ux6U_6U_1_3385_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3400
         assign bnn_Add_17Sx16S_17S_1_3400_out1 = bnn_Add_17Sx16S_17S_1_3400_in2 + {bnn_Add_17Sx16S_17S_1_3400_in1[15], bnn_Add_17Sx16S_17S_1_3400_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3387_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5003_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3401_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3401_in2 = bnn_Mod_6Ux32U_7U_4_5003_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3401_in2 = {bnn_Add_5Sx4S_6S_1_3387_out1[4], bnn_Add_5Sx4S_6S_1_3387_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1067[6:1] or bnn_N_Mux_2_2_3_1_3386_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3401_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3401_in1 = s_reg_1067[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3401_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3386_out1[1]}}, bnn_N_Mux_2_2_3_1_3386_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3401
         assign bnn_Add_6Ux6U_6U_1_3401_out1 = bnn_Add_6Ux6U_6U_1_3401_in2 + bnn_Add_6Ux6U_6U_1_3401_in1;

         // resource: mux_2bx2i
         always @(s_reg_971 or bnn_N_Mux_2_2_3_1_1990_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3402_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3402_in3 = s_reg_971;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3402_in3 = bnn_N_Mux_2_2_3_1_1990_out1;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_Minus_2S_2S_1_1409_out1 or bnn_Minus_2S_2S_1_3379_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3402_in2
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3402_in2 = bnn_Minus_2S_2S_1_1409_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3402_in2 = bnn_Minus_2S_2S_1_3379_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_3402_in3 or bnn_N_Mux_2_2_3_1_3402_in2)
          begin :bnn_N_Mux_2_2_3_1_3402
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3402_out1 = bnn_N_Mux_2_2_3_1_3402_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3402_out1 = bnn_N_Mux_2_2_3_1_3402_in3;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3403
         assign bnn_Add_5Sx4S_6S_1_3403_out1 = {bnn_Add_5Sx4S_6S_1_3390_out1[4], bnn_Add_5Sx4S_6S_1_3390_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3389_out1[1]}}, bnn_N_Mux_2_2_3_1_3389_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_3402_in3 or bnn_N_Mux_2_2_3_1_3402_in2)
          begin :bnn_N_Mux_2_2_3_1_3405
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3405_out1 = bnn_N_Mux_2_2_3_1_3402_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3405_out1 = bnn_N_Mux_2_2_3_1_3402_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1136 or bnn_Add_4Sx2S_5S_1_2315_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3406_in2
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3406_in2 = bnn_Add_4Sx2S_5S_1_2315_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3406_in2 = s_reg_1136;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_N_Mux_2_2_3_1_1406_out1 or bnn_N_Mux_2_2_3_1_3392_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3406_in1
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3406_in1_slice = bnn_N_Mux_2_2_3_1_1406_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3406_in1_slice = bnn_N_Mux_2_2_3_1_3392_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3406
         assign bnn_Add_5Sx4S_6S_1_3406_out1 = {bnn_Add_5Sx4S_6S_1_3406_in2[4], bnn_Add_5Sx4S_6S_1_3406_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_3406_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_3406_in1_slice};

         // resource: mux_2bx2i
         always @(s_reg_979 or bnn_N_Mux_2_2_3_1_2181_out1 or gs_ctrl105)
          begin :drive_bnn_Minus_2S_2S_4_3407_in1
            if (gs_ctrl105) begin
               bnn_Minus_2S_2S_4_3407_in1 = s_reg_979;
            end
            else begin
               bnn_Minus_2S_2S_4_3407_in1 = bnn_N_Mux_2_2_3_1_2181_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_4  instance: bnn_Minus_2S_2S_4_3407
         assign bnn_Minus_2S_2S_4_3407_out1 = -bnn_Minus_2S_2S_4_3407_in1;

         // resource: mux_2bx2i
         always @(s_reg_974 or bnn_N_Mux_2_2_3_1_2001_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_4_3408_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_4_3408_in3 = s_reg_974;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3408_in3 = bnn_N_Mux_2_2_3_1_2001_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_Minus_2S_2S_4_3393_out1 or bnn_N_Mux_2_2_3_4_3408_in3)
          begin :bnn_N_Mux_2_2_3_4_3408
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3408_out1 = bnn_Minus_2S_2S_4_3393_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3408_out1 = bnn_N_Mux_2_2_3_4_3408_in3;
            end
         end

         // resource: mux_5bx2i
         always @(s_reg_1130 or bnn_Add_4Sx2S_5S_1_2343_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3409_in2
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3409_in2 = bnn_Add_4Sx2S_5S_1_2343_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3409_in2 = s_reg_1130;
            end
         end

         // resource: mux_2bx2i
         always @(bnn_N_Mux_2_2_3_1_3394_out1 or bnn_N_Mux_2_2_3_1_3780_out1 or gs_ctrl105)
          begin :drive_bnn_Add_5Sx4S_6S_1_3409_in1
            if (gs_ctrl105) begin
               bnn_Add_5Sx4S_6S_1_3409_in1_slice = bnn_N_Mux_2_2_3_1_3780_out1;
            end
            else begin
               bnn_Add_5Sx4S_6S_1_3409_in1_slice = bnn_N_Mux_2_2_3_1_3394_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3409
         assign bnn_Add_5Sx4S_6S_1_3409_out1 = {bnn_Add_5Sx4S_6S_1_3409_in2[4], bnn_Add_5Sx4S_6S_1_3409_in2} + {{ 4 {bnn_Add_5Sx4S_6S_1_3409_in1_slice[1]}}, bnn_Add_5Sx4S_6S_1_3409_in1_slice};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3410
         assign bnn_Minus_2S_2S_1_3410_out1 = -bnn_N_Mux_2_2_3_1_2012_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2199_out1 or bnn_Minus_2S_2S_4_3395_out1)
          begin :bnn_N_Mux_2_2_3_4_3411
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_3411_out1 = bnn_Minus_2S_2S_4_3395_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3411_out1 = bnn_N_Mux_2_2_3_1_2199_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3412_in3 = {bnn_RightShift_64Sx8S_1S_4_3397_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3398_out1 or bnn_N_Mux_2_2_3_4_3412_in3)
          begin :bnn_N_Mux_2_2_3_4_3412
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3412_out1 = bnn_N_Mux_2_2_3_4_3398_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3412_out1 = bnn_N_Mux_2_2_3_4_3412_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3413_in1 = {s_reg_1058_stage1_slice[4:0], 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3413
         assign bnn_RightShift_64Sx8S_1S_4_3413_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3413_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3399_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3414
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3414_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3414_out1 = bnn_N_Mux_2_4_8_4_3399_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3415_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[55], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2137_out1 or bnn_N_Mux_2_2_3_1_2140_out1 or bnn_N_Mux_2_2_3_4_2146_out1 or bnn_N_Mux_2_4_8_4_3415_in3)
          begin :bnn_N_Mux_2_4_8_4_3415
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3415_out1 = bnn_N_Mux_2_2_3_1_2137_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3415_out1 = bnn_N_Mux_2_4_8_4_3415_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3415_out1 = bnn_N_Mux_2_2_3_1_2140_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3415_out1 = bnn_N_Mux_2_2_3_4_2146_out1;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2211_out1 or bnn_N_Mux_2_2_3_1_2214_out1 or bnn_N_Mux_2_4_8_4_3415_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3416
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3416_out1 = bnn_N_Mux_2_2_3_1_2211_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3416_out1 = bnn_N_Mux_2_4_8_4_3415_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3416_out1 = bnn_N_Mux_2_2_3_1_2214_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3416_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3417
         assign bnn_RightShift_64Sx8S_1S_4_3417_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_Sub_8Sx2S_8S_4_1619_out1[5:0];

         // resource: mux_17bx2i
         always @(fixed_buffer_52_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4607_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3418_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3418_in2 = {bnn_Mul_16Sx12S_19S_4_4607_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3418_in2 = {{ 5 {fixed_buffer_52_if_1_dout_wire[11]}}, fixed_buffer_52_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3401_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3418_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3418_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3418_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3401_out1[4]}}, bnn_Add_6Ux6U_6U_1_3401_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3418
         assign bnn_Add_17Sx16S_17S_1_3418_out1 = bnn_Add_17Sx16S_17S_1_3418_in2 + {bnn_Add_17Sx16S_17S_1_3418_in1[15], bnn_Add_17Sx16S_17S_1_3418_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3403_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5004_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3419_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3419_in2 = bnn_Mod_6Ux32U_7U_4_5004_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3419_in2 = {bnn_Add_5Sx4S_6S_1_3403_out1[4], bnn_Add_5Sx4S_6S_1_3403_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1058[6:1] or bnn_N_Mux_2_2_3_1_3402_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3419_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3419_in1 = s_reg_1058[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3419_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3402_out1[1]}}, bnn_N_Mux_2_2_3_1_3402_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3419
         assign bnn_Add_6Ux6U_6U_1_3419_out1 = bnn_Add_6Ux6U_6U_1_3419_in2 + bnn_Add_6Ux6U_6U_1_3419_in1;

         // resource: mux_2bx2i
         always @(bnn_Minus_2S_2S_1_1423_out1 or bnn_Minus_2S_2S_4_3393_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_1_3420_in2
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_1_3420_in2 = bnn_Minus_2S_2S_1_1423_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3420_in2 = bnn_Minus_2S_2S_4_3393_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_N_Mux_2_2_3_4_3408_in3 or bnn_N_Mux_2_2_3_1_3420_in2)
          begin :bnn_N_Mux_2_2_3_1_3420
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_3420_out1 = bnn_N_Mux_2_2_3_1_3420_in2;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3420_out1 = bnn_N_Mux_2_2_3_4_3408_in3;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3421
         assign bnn_Add_5Sx4S_6S_1_3421_out1 = {bnn_Add_5Sx4S_6S_1_3406_out1[4], bnn_Add_5Sx4S_6S_1_3406_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3405_out1[1]}}, bnn_N_Mux_2_2_3_1_3405_out1};

         // resource: mux_2bx2i
         always @(s_reg_979 or bnn_N_Mux_2_2_3_1_2181_out1 or gs_ctrl105)
          begin :drive_bnn_N_Mux_2_2_3_4_3423_in3
            if (gs_ctrl105) begin
               bnn_N_Mux_2_2_3_4_3423_in3 = s_reg_979;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3423_in3 = bnn_N_Mux_2_2_3_1_2181_out1;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_4_3407_out1 or bnn_N_Mux_2_2_3_4_3423_in3)
          begin :bnn_N_Mux_2_2_3_4_3423
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3423_out1 = bnn_Minus_2S_2S_4_3407_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3423_out1 = bnn_N_Mux_2_2_3_4_3423_in3;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3424
         assign bnn_Add_5Sx4S_6S_1_3424_out1 = {bnn_Add_5Sx4S_6S_1_3409_out1[4], bnn_Add_5Sx4S_6S_1_3409_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3408_out1[1]}}, bnn_N_Mux_2_2_3_4_3408_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3425
         assign bnn_Minus_2S_2S_1_3425_out1 = -bnn_N_Mux_2_2_3_1_2029_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2012_out1 or bnn_Minus_2S_2S_1_3410_out1)
          begin :bnn_N_Mux_2_2_3_4_3426
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3426_out1 = bnn_Minus_2S_2S_1_3410_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3426_out1 = bnn_N_Mux_2_2_3_1_2012_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_4  instance: bnn_Add_5Sx4S_6S_4_3427
         assign bnn_Add_5Sx4S_6S_4_3427_out1 = {s_reg_1137[4], s_reg_1137} + {{ 4 {bnn_N_Mux_2_2_3_4_3411_out1[1]}}, bnn_N_Mux_2_2_3_4_3411_out1};

         assign bnn_N_Mux_2_2_3_4_3428_in3 = {bnn_RightShift_64Sx8S_1S_4_3413_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3414_out1 or bnn_N_Mux_2_2_3_4_3428_in3)
          begin :bnn_N_Mux_2_2_3_4_3428
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3428_out1 = bnn_N_Mux_2_2_3_4_3414_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3428_out1 = bnn_N_Mux_2_2_3_4_3428_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3429_in1 = {s_reg_1058_stage1_slice[4:0], 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3429
         assign bnn_RightShift_64Sx8S_1S_4_3429_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3429_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3415_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3430
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3430_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3430_out1 = bnn_N_Mux_2_4_8_4_3415_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3431_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[56], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2193_out1 or bnn_N_Mux_2_2_3_1_2196_out1 or bnn_N_Mux_2_4_8_4_3431_in3 or bnn_N_Mux_3_2_6_4_1833_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3431
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3431_out1 = bnn_N_Mux_2_2_3_1_2193_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3431_out1 = bnn_N_Mux_2_4_8_4_3431_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3431_out1 = bnn_N_Mux_2_2_3_1_2196_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3431_out1 = bnn_N_Mux_3_2_6_4_1833_out1_slice;
               end
               
            endcase

         end

         assign bnn_RightShift_64Sx8S_1S_4_3432_in1 = {s_reg_1110, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3432
         assign bnn_RightShift_64Sx8S_1S_4_3432_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3432_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3416_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3433
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3433_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3433_out1 = bnn_N_Mux_2_4_8_4_3416_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_4_3434_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_4_3417_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_3434_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_3434
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_3434_out1_slice = bnn_N_Mux_3_2_6_4_3434_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_3434_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2024_out1 or bnn_N_Mux_2_2_3_1_2027_out1 or bnn_N_Mux_2_4_8_4_3431_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3435
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3435_out1 = bnn_N_Mux_2_2_3_1_2024_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3435_out1 = bnn_N_Mux_2_4_8_4_3431_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3435_out1 = bnn_N_Mux_2_2_3_1_2027_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3435_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_53_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4616_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3436_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3436_in2 = {bnn_Mul_16Sx12S_19S_4_4616_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3436_in2 = {{ 5 {fixed_buffer_53_if_1_dout_wire[11]}}, fixed_buffer_53_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3419_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3436_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3436_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3436_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3419_out1[4]}}, bnn_Add_6Ux6U_6U_1_3419_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3436
         assign bnn_Add_17Sx16S_17S_1_3436_out1 = bnn_Add_17Sx16S_17S_1_3436_in2 + {bnn_Add_17Sx16S_17S_1_3436_in1[15], bnn_Add_17Sx16S_17S_1_3436_in1};

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3421_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5005_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3437_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3437_in2 = bnn_Mod_6Ux32U_7U_4_5005_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3437_in2 = {bnn_Add_5Sx4S_6S_1_3421_out1[4], bnn_Add_5Sx4S_6S_1_3421_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1046[6:1] or bnn_N_Mux_2_2_3_1_3420_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3437_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3437_in1 = s_reg_1046[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3437_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_3420_out1[1]}}, bnn_N_Mux_2_2_3_1_3420_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3437
         assign bnn_Add_6Ux6U_6U_1_3437_out1 = bnn_Add_6Ux6U_6U_1_3437_in2 + bnn_Add_6Ux6U_6U_1_3437_in1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2012_out1 or bnn_Minus_2S_2S_1_3410_out1)
          begin :bnn_N_Mux_2_2_3_1_3439
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3439_out1 = bnn_Minus_2S_2S_1_3410_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3439_out1 = bnn_N_Mux_2_2_3_1_2012_out1;
            end
         end

         // resource: mux_6bx2i
         always @(bnn_Add_5Sx4S_6S_1_3424_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5006_out1[6:1] or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3441_in2
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3441_in2 = bnn_Mod_6Ux32U_7U_4_5006_out1[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3441_in2 = {bnn_Add_5Sx4S_6S_1_3424_out1[4], bnn_Add_5Sx4S_6S_1_3424_out1[4:0]};
            end
         end

         // resource: mux_6bx2i
         always @(s_reg_1041[6:1] or bnn_N_Mux_2_2_3_4_3423_out1 or gs_ctrl61)
          begin :drive_bnn_Add_6Ux6U_6U_1_3441_in1
            if (gs_ctrl61) begin
               bnn_Add_6Ux6U_6U_1_3441_in1 = s_reg_1041[6:1];
            end
            else begin
               bnn_Add_6Ux6U_6U_1_3441_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3423_out1[1]}}, bnn_N_Mux_2_2_3_4_3423_out1};
            end
         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3441
         assign bnn_Add_6Ux6U_6U_1_3441_out1 = bnn_Add_6Ux6U_6U_1_3441_in2 + bnn_Add_6Ux6U_6U_1_3441_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2029_out1 or bnn_Minus_2S_2S_1_3425_out1)
          begin :bnn_N_Mux_2_2_3_4_3442
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3442_out1 = bnn_Minus_2S_2S_1_3425_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3442_out1 = bnn_N_Mux_2_2_3_1_2029_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3443
         assign bnn_Add_5Sx4S_6S_1_3443_out1 = {bnn_Add_5Sx4S_6S_4_3427_out1[4], bnn_Add_5Sx4S_6S_4_3427_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3426_out1[1]}}, bnn_N_Mux_2_2_3_4_3426_out1};

         assign bnn_N_Mux_2_2_3_4_3444_in3 = {bnn_RightShift_64Sx8S_1S_4_3429_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3430_out1 or bnn_N_Mux_2_2_3_4_3444_in3)
          begin :bnn_N_Mux_2_2_3_4_3444
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3444_out1 = bnn_N_Mux_2_2_3_4_3430_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3444_out1 = bnn_N_Mux_2_2_3_4_3444_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3431_out1 or s_reg_1075_stage1)
          begin :bnn_N_Mux_2_2_3_4_3445
            if (s_reg_1075_stage1) begin
               bnn_N_Mux_2_2_3_4_3445_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3445_out1 = bnn_N_Mux_2_4_8_4_3431_out1;
            end
         end

         assign bnn_N_Mux_3_2_6_4_3446_in2 = {{ 2 {bnn_RightShift_64Sx8S_1S_4_3432_out1}}, 1'b1};

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1078 or bnn_N_Mux_3_2_6_4_3446_in2[1:0])
          begin :bnn_N_Mux_3_2_6_4_3446
            if (s_reg_1078) begin
               bnn_N_Mux_3_2_6_4_3446_out1_slice = bnn_N_Mux_3_2_6_4_3446_in2[1:0];
            end
            else begin
               bnn_N_Mux_3_2_6_4_3446_out1_slice = 2'd0;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3433_out1 or bnn_N_Mux_3_2_6_4_3434_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_3447
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3447_out1 = bnn_N_Mux_2_2_3_4_3433_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3447_out1 = bnn_N_Mux_3_2_6_4_3434_out1_slice;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3448_in1 = {s_reg_1067_stage1_slice, 3'd0};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3448
         assign bnn_RightShift_64Sx8S_1S_4_3448_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3448_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3435_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3449
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3449_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3449_out1 = bnn_N_Mux_2_4_8_4_3435_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3450_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[57], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2041_out1 or bnn_N_Mux_2_2_3_1_2044_out1 or bnn_N_Mux_2_4_8_4_3450_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3450
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3450_out1 = bnn_N_Mux_2_2_3_1_2041_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3450_out1 = bnn_N_Mux_2_4_8_4_3450_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3450_out1 = bnn_N_Mux_2_2_3_1_2044_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3450_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_54_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4625_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3451_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3451_in2 = {bnn_Mul_16Sx12S_19S_4_4625_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3451_in2 = {{ 5 {fixed_buffer_54_if_1_dout_wire[11]}}, fixed_buffer_54_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3437_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3451_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3451_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3451_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3437_out1[4]}}, bnn_Add_6Ux6U_6U_1_3437_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3451
         assign bnn_Add_17Sx16S_17S_1_3451_out1 = bnn_Add_17Sx16S_17S_1_3451_in2 + {bnn_Add_17Sx16S_17S_1_3451_in1[15], bnn_Add_17Sx16S_17S_1_3451_in1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3452
         assign bnn_Minus_2S_2S_1_3452_out1 = -bnn_N_Mux_2_2_3_1_2046_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2029_out1 or bnn_Minus_2S_2S_1_3425_out1)
          begin :bnn_N_Mux_2_2_3_4_3453
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3453_out1 = bnn_Minus_2S_2S_1_3425_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3453_out1 = bnn_N_Mux_2_2_3_1_2029_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3454
         assign bnn_Add_5Sx4S_6S_1_3454_out1 = {s_reg_1138[4], s_reg_1138[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3439_out1[1]}}, bnn_N_Mux_2_2_3_1_3439_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2029_out1 or bnn_Minus_2S_2S_1_3425_out1)
          begin :bnn_N_Mux_2_2_3_1_3456
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3456_out1 = bnn_Minus_2S_2S_1_3425_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3456_out1 = bnn_N_Mux_2_2_3_1_2029_out1;
            end
         end

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1428_out1[4:0] or bnn_Add_5Sx4S_6S_1_3443_out1[4:0] or bnn_Mod_6Ux32U_7U_4_4990_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3458_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3458_in2 = {bnn_Add_5Sx4S_6S_1_1428_out1[4], bnn_Add_5Sx4S_6S_1_1428_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3458_in2 = bnn_Mod_6Ux32U_7U_4_4990_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3458_in2 = {bnn_Add_5Sx4S_6S_1_3443_out1[4], bnn_Add_5Sx4S_6S_1_3443_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1104[6:1] or bnn_N_Mux_2_2_3_1_1427_out1 or bnn_N_Mux_2_2_3_4_3442_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3458_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3458_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1427_out1[1]}}, bnn_N_Mux_2_2_3_1_1427_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3458_in1 = s_reg_1104[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3458_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3442_out1[1]}}, bnn_N_Mux_2_2_3_4_3442_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3458
         assign bnn_Add_6Ux6U_6U_1_3458_out1 = bnn_Add_6Ux6U_6U_1_3458_in2 + bnn_Add_6Ux6U_6U_1_3458_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_Or_1Sx1U_1S_4_1588_out1 or bnn_N_Mux_2_2_3_4_3445_out1 or bnn_N_Mux_3_2_6_4_3446_out1_slice)
          begin :bnn_N_Mux_2_2_3_4_3459
            if (bnn_Or_1Sx1U_1S_4_1588_out1) begin
               bnn_N_Mux_2_2_3_4_3459_out1 = bnn_N_Mux_2_2_3_4_3445_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3459_out1 = bnn_N_Mux_3_2_6_4_3446_out1_slice;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3460_in3 = {bnn_RightShift_64Sx8S_1S_4_3448_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3449_out1 or bnn_N_Mux_2_2_3_4_3460_in3)
          begin :bnn_N_Mux_2_2_3_4_3460
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3460_out1 = bnn_N_Mux_2_2_3_4_3449_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3460_out1 = bnn_N_Mux_2_2_3_4_3460_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3461_in1 = {s_reg_1067_stage1_slice, 3'd1};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3461
         assign bnn_RightShift_64Sx8S_1S_4_3461_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3461_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3450_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3462
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3462_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3462_out1 = bnn_N_Mux_2_4_8_4_3450_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3463_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[58], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2058_out1 or bnn_N_Mux_2_2_3_1_2061_out1 or bnn_N_Mux_2_4_8_4_3463_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3463
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3463_out1 = bnn_N_Mux_2_2_3_1_2058_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3463_out1 = bnn_N_Mux_2_4_8_4_3463_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3463_out1 = bnn_N_Mux_2_2_3_1_2061_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3463_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_55_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4634_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3464_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3464_in2 = {bnn_Mul_16Sx12S_19S_4_4634_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3464_in2 = {{ 5 {fixed_buffer_55_if_1_dout_wire[11]}}, fixed_buffer_55_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3441_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3464_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3464_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3464_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3441_out1[4]}}, bnn_Add_6Ux6U_6U_1_3441_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3464
         assign bnn_Add_17Sx16S_17S_1_3464_out1 = bnn_Add_17Sx16S_17S_1_3464_in2 + {bnn_Add_17Sx16S_17S_1_3464_in1[15], bnn_Add_17Sx16S_17S_1_3464_in1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2046_out1 or bnn_Minus_2S_2S_1_3452_out1)
          begin :bnn_N_Mux_2_2_3_4_3465
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3465_out1 = bnn_Minus_2S_2S_1_3452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3465_out1 = bnn_N_Mux_2_2_3_1_2046_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3466
         assign bnn_Add_5Sx4S_6S_1_3466_out1 = {bnn_Add_5Sx4S_6S_1_3454_out1[4], bnn_Add_5Sx4S_6S_1_3454_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3453_out1[1]}}, bnn_N_Mux_2_2_3_4_3453_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3467
         assign bnn_Minus_2S_2S_1_3467_out1 = -bnn_N_Mux_2_2_3_1_2063_out1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2046_out1 or bnn_Minus_2S_2S_1_3452_out1)
          begin :bnn_N_Mux_2_2_3_4_3468
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3468_out1 = bnn_Minus_2S_2S_1_3452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3468_out1 = bnn_N_Mux_2_2_3_1_2046_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3469
         assign bnn_Add_5Sx4S_6S_1_3469_out1 = {s_reg_1139[4], s_reg_1139} + {{ 4 {bnn_N_Mux_2_2_3_1_3456_out1[1]}}, bnn_N_Mux_2_2_3_1_3456_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2046_out1 or bnn_Minus_2S_2S_1_3452_out1)
          begin :bnn_N_Mux_2_2_3_1_3471
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3471_out1 = bnn_Minus_2S_2S_1_3452_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3471_out1 = bnn_N_Mux_2_2_3_1_2046_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3473_in3 = {bnn_RightShift_64Sx8S_1S_4_3461_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3462_out1 or bnn_N_Mux_2_2_3_4_3473_in3)
          begin :bnn_N_Mux_2_2_3_4_3473
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3473_out1 = bnn_N_Mux_2_2_3_4_3462_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3473_out1 = bnn_N_Mux_2_2_3_4_3473_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3474_in1 = {s_reg_1067_stage1_slice, 3'd2};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3474
         assign bnn_RightShift_64Sx8S_1S_4_3474_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3474_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3463_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3475
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3475_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3475_out1 = bnn_N_Mux_2_4_8_4_3463_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3476_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[59], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2075_out1 or bnn_N_Mux_2_2_3_1_2078_out1 or bnn_N_Mux_2_4_8_4_3476_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3476
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3476_out1 = bnn_N_Mux_2_2_3_1_2075_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3476_out1 = bnn_N_Mux_2_4_8_4_3476_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3476_out1 = bnn_N_Mux_2_2_3_1_2078_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3476_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_56_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4643_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3477_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3477_in2 = {bnn_Mul_16Sx12S_19S_4_4643_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3477_in2 = {{ 5 {fixed_buffer_56_if_1_dout_wire[11]}}, fixed_buffer_56_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3458_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3477_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3477_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3477_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3458_out1[4]}}, bnn_Add_6Ux6U_6U_1_3458_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3477
         assign bnn_Add_17Sx16S_17S_1_3477_out1 = bnn_Add_17Sx16S_17S_1_3477_in2 + {bnn_Add_17Sx16S_17S_1_3477_in1[15], bnn_Add_17Sx16S_17S_1_3477_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1445_out1[4:0] or bnn_Add_5Sx4S_6S_1_3466_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5007_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3478_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3478_in2 = {bnn_Add_5Sx4S_6S_1_1445_out1[4], bnn_Add_5Sx4S_6S_1_1445_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3478_in2 = bnn_Mod_6Ux32U_7U_4_5007_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3478_in2 = {bnn_Add_5Sx4S_6S_1_3466_out1[4], bnn_Add_5Sx4S_6S_1_3466_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1034[6:1] or bnn_N_Mux_2_2_3_1_1444_out1 or bnn_N_Mux_2_2_3_4_3465_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3478_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3478_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1444_out1[1]}}, bnn_N_Mux_2_2_3_1_1444_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3478_in1 = s_reg_1034[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3478_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3465_out1[1]}}, bnn_N_Mux_2_2_3_4_3465_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3478
         assign bnn_Add_6Ux6U_6U_1_3478_out1 = bnn_Add_6Ux6U_6U_1_3478_in2 + bnn_Add_6Ux6U_6U_1_3478_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2063_out1 or bnn_Minus_2S_2S_1_3467_out1)
          begin :bnn_N_Mux_2_2_3_4_3479
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3479_out1 = bnn_Minus_2S_2S_1_3467_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3479_out1 = bnn_N_Mux_2_2_3_1_2063_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3480
         assign bnn_Add_5Sx4S_6S_1_3480_out1 = {bnn_Add_5Sx4S_6S_1_3469_out1[4], bnn_Add_5Sx4S_6S_1_3469_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_4_3468_out1[1]}}, bnn_N_Mux_2_2_3_4_3468_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3481
         assign bnn_Minus_2S_2S_1_3481_out1 = -bnn_N_Mux_2_2_3_1_2080_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2063_out1 or bnn_Minus_2S_2S_1_3467_out1)
          begin :bnn_N_Mux_2_2_3_1_3482
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3482_out1 = bnn_Minus_2S_2S_1_3467_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3482_out1 = bnn_N_Mux_2_2_3_1_2063_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3483
         assign bnn_Add_5Sx4S_6S_1_3483_out1 = {s_reg_1140[4], s_reg_1140} + {{ 4 {bnn_N_Mux_2_2_3_1_3471_out1[1]}}, bnn_N_Mux_2_2_3_1_3471_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2063_out1 or bnn_Minus_2S_2S_1_3467_out1)
          begin :bnn_N_Mux_2_2_3_1_3485
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3485_out1 = bnn_Minus_2S_2S_1_3467_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3485_out1 = bnn_N_Mux_2_2_3_1_2063_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3487_in3 = {bnn_RightShift_64Sx8S_1S_4_3474_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3475_out1 or bnn_N_Mux_2_2_3_4_3487_in3)
          begin :bnn_N_Mux_2_2_3_4_3487
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3487_out1 = bnn_N_Mux_2_2_3_4_3475_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3487_out1 = bnn_N_Mux_2_2_3_4_3487_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3488_in1 = {s_reg_1067_stage1_slice, 3'd3};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3488
         assign bnn_RightShift_64Sx8S_1S_4_3488_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3488_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3476_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3489
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3489_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3489_out1 = bnn_N_Mux_2_4_8_4_3476_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3490_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[60], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2092_out1 or bnn_N_Mux_2_2_3_1_2095_out1 or bnn_N_Mux_2_4_8_4_3490_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3490
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3490_out1 = bnn_N_Mux_2_2_3_1_2092_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3490_out1 = bnn_N_Mux_2_4_8_4_3490_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3490_out1 = bnn_N_Mux_2_2_3_1_2095_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3490_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_57_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4652_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3491_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3491_in2 = {bnn_Mul_16Sx12S_19S_4_4652_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3491_in2 = {{ 5 {fixed_buffer_57_if_1_dout_wire[11]}}, fixed_buffer_57_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3478_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3491_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3491_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3491_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3478_out1[4]}}, bnn_Add_6Ux6U_6U_1_3478_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3491
         assign bnn_Add_17Sx16S_17S_1_3491_out1 = bnn_Add_17Sx16S_17S_1_3491_in2 + {bnn_Add_17Sx16S_17S_1_3491_in1[15], bnn_Add_17Sx16S_17S_1_3491_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1462_out1[4:0] or bnn_Add_5Sx4S_6S_1_3480_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5008_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3492_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3492_in2 = {bnn_Add_5Sx4S_6S_1_1462_out1[4], bnn_Add_5Sx4S_6S_1_1462_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3492_in2 = bnn_Mod_6Ux32U_7U_4_5008_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3492_in2 = {bnn_Add_5Sx4S_6S_1_3480_out1[4], bnn_Add_5Sx4S_6S_1_3480_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1020[6:1] or bnn_N_Mux_2_2_3_1_1461_out1 or bnn_N_Mux_2_2_3_4_3479_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3492_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3492_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1461_out1[1]}}, bnn_N_Mux_2_2_3_1_1461_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3492_in1 = s_reg_1020[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3492_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3479_out1[1]}}, bnn_N_Mux_2_2_3_4_3479_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3492
         assign bnn_Add_6Ux6U_6U_1_3492_out1 = bnn_Add_6Ux6U_6U_1_3492_in2 + bnn_Add_6Ux6U_6U_1_3492_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2080_out1 or bnn_Minus_2S_2S_1_3481_out1)
          begin :bnn_N_Mux_2_2_3_4_3493
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3493_out1 = bnn_Minus_2S_2S_1_3481_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3493_out1 = bnn_N_Mux_2_2_3_1_2080_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3494
         assign bnn_Add_5Sx4S_6S_1_3494_out1 = {bnn_Add_5Sx4S_6S_1_3483_out1[4], bnn_Add_5Sx4S_6S_1_3483_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3482_out1[1]}}, bnn_N_Mux_2_2_3_1_3482_out1};

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3495
         assign bnn_Minus_2S_2S_1_3495_out1 = -bnn_N_Mux_2_2_3_1_2097_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2080_out1 or bnn_Minus_2S_2S_1_3481_out1)
          begin :bnn_N_Mux_2_2_3_1_3496
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3496_out1 = bnn_Minus_2S_2S_1_3481_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3496_out1 = bnn_N_Mux_2_2_3_1_2080_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3497
         assign bnn_Add_5Sx4S_6S_1_3497_out1 = {s_reg_1141[4], s_reg_1141} + {{ 4 {bnn_N_Mux_2_2_3_1_3485_out1[1]}}, bnn_N_Mux_2_2_3_1_3485_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2080_out1 or bnn_Minus_2S_2S_1_3481_out1)
          begin :bnn_N_Mux_2_2_3_1_3499
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3499_out1 = bnn_Minus_2S_2S_1_3481_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3499_out1 = bnn_N_Mux_2_2_3_1_2080_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3501
         assign bnn_Minus_2S_2S_1_3501_out1 = -bnn_N_Mux_2_2_3_1_2114_out1;

         assign bnn_N_Mux_2_2_3_4_3502_in3 = {bnn_RightShift_64Sx8S_1S_4_3488_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3489_out1 or bnn_N_Mux_2_2_3_4_3502_in3)
          begin :bnn_N_Mux_2_2_3_4_3502
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3502_out1 = bnn_N_Mux_2_2_3_4_3489_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3502_out1 = bnn_N_Mux_2_2_3_4_3502_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3503_in1 = {s_reg_1067_stage1_slice, 3'd4};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3503
         assign bnn_RightShift_64Sx8S_1S_4_3503_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3503_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3490_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3504
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3504_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3504_out1 = bnn_N_Mux_2_4_8_4_3490_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3505_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[61], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2109_out1 or bnn_N_Mux_2_2_3_1_2112_out1 or bnn_N_Mux_2_4_8_4_3505_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3505
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3505_out1 = bnn_N_Mux_2_2_3_1_2109_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3505_out1 = bnn_N_Mux_2_4_8_4_3505_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3505_out1 = bnn_N_Mux_2_2_3_1_2112_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3505_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_58_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4661_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3506_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3506_in2 = {bnn_Mul_16Sx12S_19S_4_4661_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3506_in2 = {{ 5 {fixed_buffer_58_if_1_dout_wire[11]}}, fixed_buffer_58_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3492_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3506_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3506_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3506_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3492_out1[4]}}, bnn_Add_6Ux6U_6U_1_3492_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3506
         assign bnn_Add_17Sx16S_17S_1_3506_out1 = bnn_Add_17Sx16S_17S_1_3506_in2 + {bnn_Add_17Sx16S_17S_1_3506_in1[15], bnn_Add_17Sx16S_17S_1_3506_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1477_out1[4:0] or bnn_Add_5Sx4S_6S_1_3494_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5009_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3507_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3507_in2 = {bnn_Add_5Sx4S_6S_1_1477_out1[4], bnn_Add_5Sx4S_6S_1_1477_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3507_in2 = bnn_Mod_6Ux32U_7U_4_5009_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3507_in2 = {bnn_Add_5Sx4S_6S_1_3494_out1[4], bnn_Add_5Sx4S_6S_1_3494_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1019[6:1] or bnn_N_Mux_2_2_3_1_1476_out1 or bnn_N_Mux_2_2_3_4_3493_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3507_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3507_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1476_out1[1]}}, bnn_N_Mux_2_2_3_1_1476_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3507_in1 = s_reg_1019[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3507_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3493_out1[1]}}, bnn_N_Mux_2_2_3_4_3493_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3507
         assign bnn_Add_6Ux6U_6U_1_3507_out1 = bnn_Add_6Ux6U_6U_1_3507_in2 + bnn_Add_6Ux6U_6U_1_3507_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2097_out1 or bnn_Minus_2S_2S_1_3495_out1)
          begin :bnn_N_Mux_2_2_3_4_3508
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3508_out1 = bnn_Minus_2S_2S_1_3495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3508_out1 = bnn_N_Mux_2_2_3_1_2097_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3509
         assign bnn_Add_5Sx4S_6S_1_3509_out1 = {bnn_Add_5Sx4S_6S_1_3497_out1[4], bnn_Add_5Sx4S_6S_1_3497_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3496_out1[1]}}, bnn_N_Mux_2_2_3_1_3496_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2097_out1 or bnn_Minus_2S_2S_1_3495_out1)
          begin :bnn_N_Mux_2_2_3_1_3511
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3511_out1 = bnn_Minus_2S_2S_1_3495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3511_out1 = bnn_N_Mux_2_2_3_1_2097_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3512
         assign bnn_Add_5Sx4S_6S_1_3512_out1 = {s_reg_1142[4], s_reg_1142} + {{ 4 {bnn_N_Mux_2_2_3_1_3499_out1[1]}}, bnn_N_Mux_2_2_3_1_3499_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2097_out1 or bnn_Minus_2S_2S_1_3495_out1)
          begin :bnn_N_Mux_2_2_3_1_3514
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3514_out1 = bnn_Minus_2S_2S_1_3495_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3514_out1 = bnn_N_Mux_2_2_3_1_2097_out1;
            end
         end

         // resource: bnn_Minus_2S_2S_1  instance: bnn_Minus_2S_2S_1_3515
         assign bnn_Minus_2S_2S_1_3515_out1 = -bnn_N_Mux_2_2_3_1_2131_out1;

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_N_Mux_2_2_3_1_2114_out1 or bnn_Minus_2S_2S_1_3501_out1)
          begin :bnn_N_Mux_2_2_3_1_3516
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3516_out1 = bnn_Minus_2S_2S_1_3501_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3516_out1 = bnn_N_Mux_2_2_3_1_2114_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3517_in3 = {bnn_RightShift_64Sx8S_1S_4_3503_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3504_out1 or bnn_N_Mux_2_2_3_4_3517_in3)
          begin :bnn_N_Mux_2_2_3_4_3517
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3517_out1 = bnn_N_Mux_2_2_3_4_3504_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3517_out1 = bnn_N_Mux_2_2_3_4_3517_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3518_in1 = {s_reg_1067_stage1_slice, 3'd5};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3518
         assign bnn_RightShift_64Sx8S_1S_4_3518_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3518_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3505_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3519
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3519_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3519_out1 = bnn_N_Mux_2_4_8_4_3505_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3520_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[62], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_1_2126_out1 or bnn_N_Mux_2_2_3_1_2129_out1 or bnn_N_Mux_2_4_8_4_3520_in3 or bnn_N_Mux_3_2_6_1_1785_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3520
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3520_out1 = bnn_N_Mux_2_2_3_1_2126_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3520_out1 = bnn_N_Mux_2_4_8_4_3520_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3520_out1 = bnn_N_Mux_2_2_3_1_2129_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3520_out1 = bnn_N_Mux_3_2_6_1_1785_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_59_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4670_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3521_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3521_in2 = {bnn_Mul_16Sx12S_19S_4_4670_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3521_in2 = {{ 5 {fixed_buffer_59_if_1_dout_wire[11]}}, fixed_buffer_59_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3507_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3521_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3521_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3521_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3507_out1[4]}}, bnn_Add_6Ux6U_6U_1_3507_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3521
         assign bnn_Add_17Sx16S_17S_1_3521_out1 = bnn_Add_17Sx16S_17S_1_3521_in2 + {bnn_Add_17Sx16S_17S_1_3521_in1[15], bnn_Add_17Sx16S_17S_1_3521_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1489_out1[4:0] or bnn_Add_5Sx4S_6S_1_3509_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5010_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3522_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3522_in2 = {bnn_Add_5Sx4S_6S_1_1489_out1[4], bnn_Add_5Sx4S_6S_1_1489_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3522_in2 = bnn_Mod_6Ux32U_7U_4_5010_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3522_in2 = {bnn_Add_5Sx4S_6S_1_3509_out1[4], bnn_Add_5Sx4S_6S_1_3509_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1098[6:1] or bnn_N_Mux_2_2_3_1_1488_out1 or bnn_N_Mux_2_2_3_4_3508_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3522_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3522_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1488_out1[1]}}, bnn_N_Mux_2_2_3_1_1488_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3522_in1 = s_reg_1098[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3522_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3508_out1[1]}}, bnn_N_Mux_2_2_3_4_3508_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3522
         assign bnn_Add_6Ux6U_6U_1_3522_out1 = bnn_Add_6Ux6U_6U_1_3522_in2 + bnn_Add_6Ux6U_6U_1_3522_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2114_out1 or bnn_Minus_2S_2S_1_3501_out1)
          begin :bnn_N_Mux_2_2_3_4_3523
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3523_out1 = bnn_Minus_2S_2S_1_3501_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3523_out1 = bnn_N_Mux_2_2_3_1_2114_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3524
         assign bnn_Add_5Sx4S_6S_1_3524_out1 = {bnn_Add_5Sx4S_6S_1_3512_out1[4], bnn_Add_5Sx4S_6S_1_3512_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3511_out1[1]}}, bnn_N_Mux_2_2_3_1_3511_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2114_out1 or bnn_Minus_2S_2S_1_3501_out1)
          begin :bnn_N_Mux_2_2_3_1_3526
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3526_out1 = bnn_Minus_2S_2S_1_3501_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3526_out1 = bnn_N_Mux_2_2_3_1_2114_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3527
         assign bnn_Add_5Sx4S_6S_1_3527_out1 = {s_reg_1143[4], s_reg_1143} + {{ 4 {bnn_N_Mux_2_2_3_1_3514_out1[1]}}, bnn_N_Mux_2_2_3_1_3514_out1};

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_N_Mux_2_2_3_1_2131_out1 or bnn_Minus_2S_2S_1_3515_out1)
          begin :bnn_N_Mux_2_2_3_1_3528
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_3528_out1 = bnn_Minus_2S_2S_1_3515_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3528_out1 = bnn_N_Mux_2_2_3_1_2131_out1;
            end
         end

         assign bnn_N_Mux_2_2_3_4_3530_in3 = {bnn_RightShift_64Sx8S_1S_4_3518_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3519_out1 or bnn_N_Mux_2_2_3_4_3530_in3)
          begin :bnn_N_Mux_2_2_3_4_3530
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3530_out1 = bnn_N_Mux_2_2_3_4_3519_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3530_out1 = bnn_N_Mux_2_2_3_4_3530_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3531_in1 = {s_reg_1067_stage1_slice, 3'd6};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3531
         assign bnn_RightShift_64Sx8S_1S_4_3531_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3531_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3520_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3532
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3532_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3532_out1 = bnn_N_Mux_2_4_8_4_3520_out1;
            end
         end

         assign bnn_N_Mux_2_4_8_4_3533_in3 = {bnn_N_Mux_64_2_2_1_1636_out1[63], 1'b1};

         // resource: bnn_N_Mux_2_4_8_4
         always @(s_reg_1004 or bnn_N_Mux_2_2_3_4_2143_out1 or bnn_N_Mux_2_2_3_4_2146_out1 or bnn_N_Mux_2_4_8_4_3533_in3 or bnn_N_Mux_3_2_6_4_1922_out1_slice)
          begin :bnn_N_Mux_2_4_8_4_3533
            case (s_reg_1004) 

               2'd1: begin
                  bnn_N_Mux_2_4_8_4_3533_out1 = bnn_N_Mux_2_2_3_4_2143_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_4_8_4_3533_out1 = bnn_N_Mux_2_4_8_4_3533_in3;
               end
               
               2'd3: begin
                  bnn_N_Mux_2_4_8_4_3533_out1 = bnn_N_Mux_2_2_3_4_2146_out1;
               end
               
               default: begin
                  bnn_N_Mux_2_4_8_4_3533_out1 = bnn_N_Mux_3_2_6_4_1922_out1_slice;
               end
               
            endcase

         end

         // resource: mux_17bx2i
         always @(fixed_buffer_60_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4679_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3534_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3534_in2 = {bnn_Mul_16Sx12S_19S_4_4679_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3534_in2 = {{ 5 {fixed_buffer_60_if_1_dout_wire[11]}}, fixed_buffer_60_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3522_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3534_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3534_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3534_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3522_out1[4]}}, bnn_Add_6Ux6U_6U_1_3522_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3534
         assign bnn_Add_17Sx16S_17S_1_3534_out1 = bnn_Add_17Sx16S_17S_1_3534_in2 + {bnn_Add_17Sx16S_17S_1_3534_in1[15], bnn_Add_17Sx16S_17S_1_3534_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1389_out1[4:0] or bnn_Add_5Sx4S_6S_1_3524_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5011_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3535_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3535_in2 = {bnn_Add_5Sx4S_6S_1_1389_out1[4], bnn_Add_5Sx4S_6S_1_1389_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3535_in2 = bnn_Mod_6Ux32U_7U_4_5011_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3535_in2 = {bnn_Add_5Sx4S_6S_1_3524_out1[4], bnn_Add_5Sx4S_6S_1_3524_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1096[6:1] or bnn_N_Mux_2_2_3_1_976_out1 or bnn_N_Mux_2_2_3_4_3523_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3535_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3535_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_976_out1[1]}}, bnn_N_Mux_2_2_3_1_976_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3535_in1 = s_reg_1096[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3535_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3523_out1[1]}}, bnn_N_Mux_2_2_3_4_3523_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3535
         assign bnn_Add_6Ux6U_6U_1_3535_out1 = bnn_Add_6Ux6U_6U_1_3535_in2 + bnn_Add_6Ux6U_6U_1_3535_in1;

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_N_Mux_2_2_3_1_2131_out1 or bnn_Minus_2S_2S_1_3515_out1)
          begin :bnn_N_Mux_2_2_3_4_3536
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3536_out1 = bnn_Minus_2S_2S_1_3515_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3536_out1 = bnn_N_Mux_2_2_3_1_2131_out1;
            end
         end

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3537
         assign bnn_Add_5Sx4S_6S_1_3537_out1 = {bnn_Add_5Sx4S_6S_1_3527_out1[4], bnn_Add_5Sx4S_6S_1_3527_out1[4:0]} + {{ 4 {bnn_N_Mux_2_2_3_1_3526_out1[1]}}, bnn_N_Mux_2_2_3_1_3526_out1};

         // resource: bnn_Add_5Sx4S_6S_1  instance: bnn_Add_5Sx4S_6S_1_3538
         assign bnn_Add_5Sx4S_6S_1_3538_out1 = {bnn_Add_5Sx3S_5S_1_211_out1[4], bnn_Add_5Sx3S_5S_1_211_out1} + {{ 4 {bnn_N_Mux_2_2_3_1_3528_out1[1]}}, bnn_N_Mux_2_2_3_1_3528_out1};

         assign bnn_N_Mux_2_2_3_4_3539_in3 = {bnn_RightShift_64Sx8S_1S_4_3531_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3532_out1 or bnn_N_Mux_2_2_3_4_3539_in3)
          begin :bnn_N_Mux_2_2_3_4_3539
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3539_out1 = bnn_N_Mux_2_2_3_4_3532_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3539_out1 = bnn_N_Mux_2_2_3_4_3539_in3;
            end
         end

         assign bnn_RightShift_64Sx8S_1S_4_3540_in1 = {s_reg_1067_stage1_slice, 3'd7};

         // resource: bnn_RightShift_64Sx8S_1S_4  instance: bnn_RightShift_64Sx8S_1S_4_3540
         assign bnn_RightShift_64Sx8S_1S_4_3540_out1 = {{ 64 {bnn_N_Mux_64_2_2_1_1636_out1[63]}}, bnn_N_Mux_64_2_2_1_1636_out1} >> bnn_RightShift_64Sx8S_1S_4_3540_in1[5:0];

         // resource: bnn_N_Mux_2_2_3_4
         always @(bnn_N_Mux_2_4_8_4_3533_out1 or s_reg_1083_stage1)
          begin :bnn_N_Mux_2_2_3_4_3541
            if (s_reg_1083_stage1) begin
               bnn_N_Mux_2_2_3_4_3541_out1 = 2'd0;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3541_out1 = bnn_N_Mux_2_4_8_4_3533_out1;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_61_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4688_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3542_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3542_in2 = {bnn_Mul_16Sx12S_19S_4_4688_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3542_in2 = {{ 5 {fixed_buffer_61_if_1_dout_wire[11]}}, fixed_buffer_61_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3535_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3542_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3542_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3542_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3535_out1[4]}}, bnn_Add_6Ux6U_6U_1_3535_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3542
         assign bnn_Add_17Sx16S_17S_1_3542_out1 = bnn_Add_17Sx16S_17S_1_3542_in2 + {bnn_Add_17Sx16S_17S_1_3542_in1[15], bnn_Add_17Sx16S_17S_1_3542_in1};

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1400_out1[4:0] or bnn_Add_5Sx4S_6S_1_3537_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5012_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3543_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3543_in2 = {bnn_Add_5Sx4S_6S_1_1400_out1[4], bnn_Add_5Sx4S_6S_1_1400_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3543_in2 = bnn_Mod_6Ux32U_7U_4_5012_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3543_in2 = {bnn_Add_5Sx4S_6S_1_3537_out1[4], bnn_Add_5Sx4S_6S_1_3537_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1105[6:1] or bnn_N_Mux_2_2_3_1_1028_out1 or bnn_N_Mux_2_2_3_4_3536_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3543_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3543_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1028_out1[1]}}, bnn_N_Mux_2_2_3_1_1028_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3543_in1 = s_reg_1105[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3543_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_3536_out1[1]}}, bnn_N_Mux_2_2_3_4_3536_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3543
         assign bnn_Add_6Ux6U_6U_1_3543_out1 = bnn_Add_6Ux6U_6U_1_3543_in2 + bnn_Add_6Ux6U_6U_1_3543_in1;

         // resource: mux_6bx3i
         always @(bnn_Add_5Sx4S_6S_1_1315_out1[4:0] or bnn_Add_5Sx4S_6S_1_3538_out1[4:0] or bnn_Mod_6Ux32U_7U_4_5018_out1[6:1] or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3544_in2
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3544_in2 = {bnn_Add_5Sx4S_6S_1_1315_out1[4], bnn_Add_5Sx4S_6S_1_1315_out1[4:0]};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3544_in2 = bnn_Mod_6Ux32U_7U_4_5018_out1[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3544_in2 = {bnn_Add_5Sx4S_6S_1_3538_out1[4], bnn_Add_5Sx4S_6S_1_3538_out1[4:0]};
               end
               
            endcase

         end

         // resource: mux_6bx3i
         always @(s_reg_1086[6:1] or bnn_N_Mux_2_2_3_1_1048_out1 or bnn_N_Mux_2_2_3_4_1635_out1 or gs_ctrl23)
          begin :drive_bnn_Add_6Ux6U_6U_1_3544_in1
            case (gs_ctrl23) 

               2'd1: begin
                  bnn_Add_6Ux6U_6U_1_3544_in1 = {{ 4 {bnn_N_Mux_2_2_3_1_1048_out1[1]}}, bnn_N_Mux_2_2_3_1_1048_out1};
               end
               
               2'd2: begin
                  bnn_Add_6Ux6U_6U_1_3544_in1 = s_reg_1086[6:1];
               end
               
               default: begin
                  bnn_Add_6Ux6U_6U_1_3544_in1 = {{ 4 {bnn_N_Mux_2_2_3_4_1635_out1[1]}}, bnn_N_Mux_2_2_3_4_1635_out1};
               end
               
            endcase

         end

         // resource: bnn_Add_6Ux6U_6U_1  instance: bnn_Add_6Ux6U_6U_1_3544
         assign bnn_Add_6Ux6U_6U_1_3544_out1 = bnn_Add_6Ux6U_6U_1_3544_in2 + bnn_Add_6Ux6U_6U_1_3544_in1;

         assign bnn_N_Mux_2_2_3_4_3545_in3 = {bnn_RightShift_64Sx8S_1S_4_3540_out1, 1'b1};

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_1082 or bnn_N_Mux_2_2_3_4_3541_out1 or bnn_N_Mux_2_2_3_4_3545_in3)
          begin :bnn_N_Mux_2_2_3_4_3545
            if (s_reg_1082) begin
               bnn_N_Mux_2_2_3_4_3545_out1 = bnn_N_Mux_2_2_3_4_3541_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3545_out1 = bnn_N_Mux_2_2_3_4_3545_in3;
            end
         end

         // resource: mux_17bx2i
         always @(fixed_buffer_62_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4697_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3546_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3546_in2 = {bnn_Mul_16Sx12S_19S_4_4697_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3546_in2 = {{ 5 {fixed_buffer_62_if_1_dout_wire[11]}}, fixed_buffer_62_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3543_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3546_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3546_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3546_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3543_out1[4]}}, bnn_Add_6Ux6U_6U_1_3543_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3546
         assign bnn_Add_17Sx16S_17S_1_3546_out1 = bnn_Add_17Sx16S_17S_1_3546_in2 + {bnn_Add_17Sx16S_17S_1_3546_in1[15], bnn_Add_17Sx16S_17S_1_3546_in1};

         // resource: mux_17bx2i
         always @(fixed_buffer_63_if_1_dout_wire or bnn_Mul_16Sx12S_19S_4_4706_out1[18:3] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3547_in2
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3547_in2 = {bnn_Mul_16Sx12S_19S_4_4706_out1[18:3], 1'b0};
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3547_in2 = {{ 5 {fixed_buffer_63_if_1_dout_wire[11]}}, fixed_buffer_63_if_1_dout_wire};
            end
         end

         // resource: mux_16bx2i
         always @(s_reg_1138 or bnn_Add_6Ux6U_6U_1_3544_out1[4:0] or gs_ctrl0)
          begin :drive_bnn_Add_17Sx16S_17S_1_3547_in1
            if (gs_ctrl0) begin
               bnn_Add_17Sx16S_17S_1_3547_in1 = s_reg_1138;
            end
            else begin
               bnn_Add_17Sx16S_17S_1_3547_in1 = {{ 11 {bnn_Add_6Ux6U_6U_1_3544_out1[4]}}, bnn_Add_6Ux6U_6U_1_3544_out1[4:0]};
            end
         end

         // resource: bnn_Add_17Sx16S_17S_1  instance: bnn_Add_17Sx16S_17S_1_3547
         assign bnn_Add_17Sx16S_17S_1_3547_out1 = bnn_Add_17Sx16S_17S_1_3547_in2 + {bnn_Add_17Sx16S_17S_1_3547_in1[15], bnn_Add_17Sx16S_17S_1_3547_in1};

         // resource: bnn_OrReduction_2U_1U_4  instance: bnn_OrReduction_2U_1U_4_3548
         assign bnn_OrReduction_2U_1U_4_3548_out1 = |s_reg_1004;

         // resource: mux_2bx3i
         always @(s_reg_872 or s_reg_992 or bnn_N_Mux_2_2_3_1_3071_out1 or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_3630_in3
            case (gs_ctrl196) 

               2'd1: begin
                  bnn_N_Mux_2_2_3_1_3630_in3 = bnn_N_Mux_2_2_3_1_3071_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_3630_in3 = s_reg_992;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_3630_in3 = s_reg_872;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_1302_out1 or bnn_N_Mux_2_2_3_1_3630_in3)
          begin :bnn_N_Mux_2_2_3_1_3630
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3630_out1 = bnn_Minus_2S_2S_1_1302_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3630_out1 = bnn_N_Mux_2_2_3_1_3630_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_890 or bnn_N_Mux_2_2_3_1_3151_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_3724_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_3724_in3 = bnn_N_Mux_2_2_3_1_3151_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3724_in3 = s_reg_890;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_1_1490_out1 or bnn_N_Mux_2_2_3_4_3724_in3)
          begin :bnn_N_Mux_2_2_3_4_3724
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3724_out1 = bnn_Minus_2S_2S_1_1490_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3724_out1 = bnn_N_Mux_2_2_3_4_3724_in3;
            end
         end

         // resource: mux_2bx3i
         always @(s_reg_890 or s_reg_965 or bnn_N_Mux_2_2_3_1_3151_out1 or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_3730_in3
            case (gs_ctrl196) 

               2'd1: begin
                  bnn_N_Mux_2_2_3_1_3730_in3 = bnn_N_Mux_2_2_3_1_3151_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_3730_in3 = s_reg_965;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_3730_in3 = s_reg_890;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_1490_out1 or bnn_N_Mux_2_2_3_1_3730_in3)
          begin :bnn_N_Mux_2_2_3_1_3730
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3730_out1 = bnn_Minus_2S_2S_1_1490_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3730_out1 = bnn_N_Mux_2_2_3_1_3730_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_911 or bnn_N_Mux_2_2_3_1_3184_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_3774_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_3774_in3 = bnn_N_Mux_2_2_3_1_3184_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3774_in3 = s_reg_911;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_1_1287_out1 or bnn_N_Mux_2_2_3_4_3774_in3)
          begin :bnn_N_Mux_2_2_3_4_3774
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3774_out1 = bnn_Minus_2S_2S_1_1287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3774_out1 = bnn_N_Mux_2_2_3_4_3774_in3;
            end
         end

         // resource: mux_2bx3i
         always @(s_reg_911 or s_reg_971 or bnn_N_Mux_2_2_3_1_3184_out1 or gs_ctrl196)
          begin :drive_bnn_N_Mux_2_2_3_1_3780_in3
            case (gs_ctrl196) 

               2'd1: begin
                  bnn_N_Mux_2_2_3_1_3780_in3 = bnn_N_Mux_2_2_3_1_3184_out1;
               end
               
               2'd2: begin
                  bnn_N_Mux_2_2_3_1_3780_in3 = s_reg_971;
               end
               
               default: begin
                  bnn_N_Mux_2_2_3_1_3780_in3 = s_reg_911;
               end
               
            endcase

         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_1287_out1 or bnn_N_Mux_2_2_3_1_3780_in3)
          begin :bnn_N_Mux_2_2_3_1_3780
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_3780_out1 = bnn_Minus_2S_2S_1_1287_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_3780_out1 = bnn_N_Mux_2_2_3_1_3780_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_886[1:0] or bnn_N_Mux_2_2_3_1_3216_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_3827_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_3827_in3 = bnn_N_Mux_2_2_3_1_3216_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3827_in3 = s_reg_886[1:0];
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_Minus_2S_2S_1_1299_out1 or bnn_N_Mux_2_2_3_4_3827_in3)
          begin :bnn_N_Mux_2_2_3_4_3827
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_3827_out1 = bnn_Minus_2S_2S_1_1299_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3827_out1 = bnn_N_Mux_2_2_3_4_3827_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_895 or bnn_N_Mux_2_2_3_1_3229_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_3849_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_3849_in3 = bnn_N_Mux_2_2_3_1_3229_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3849_in3 = s_reg_895;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_1_1392_out1 or bnn_N_Mux_2_2_3_4_3849_in3)
          begin :bnn_N_Mux_2_2_3_4_3849
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_3849_out1 = bnn_Minus_2S_2S_1_1392_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_3849_out1 = bnn_N_Mux_2_2_3_4_3849_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_943 or bnn_N_Mux_2_2_3_4_3325_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_4010_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_1_4010_in3 = bnn_N_Mux_2_2_3_4_3325_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4010_in3 = s_reg_943;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_1503_out1 or bnn_N_Mux_2_2_3_1_4010_in3)
          begin :bnn_N_Mux_2_2_3_1_4010
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_4010_out1 = bnn_Minus_2S_2S_1_1503_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4010_out1 = bnn_N_Mux_2_2_3_1_4010_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_949 or bnn_N_Mux_2_2_3_1_3338_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_4032_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_4032_in3 = bnn_N_Mux_2_2_3_1_3338_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4032_in3 = s_reg_949;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_Minus_2S_2S_1_1404_out1 or bnn_N_Mux_2_2_3_4_4032_in3)
          begin :bnn_N_Mux_2_2_3_4_4032
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_4032_out1 = bnn_Minus_2S_2S_1_1404_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4032_out1 = bnn_N_Mux_2_2_3_4_4032_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_955 or bnn_N_Mux_2_2_3_4_3351_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_4_4054_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_4_4054_in3 = bnn_N_Mux_2_2_3_4_3351_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4054_in3 = s_reg_955;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_957 or bnn_Minus_2S_2S_4_960_out1 or bnn_N_Mux_2_2_3_4_4054_in3)
          begin :bnn_N_Mux_2_2_3_4_4054
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_4_4054_out1 = bnn_Minus_2S_2S_4_960_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4054_out1 = bnn_N_Mux_2_2_3_4_4054_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_951 or bnn_Minus_2S_2S_4_960_out1 or bnn_N_Mux_2_2_3_4_4054_in3)
          begin :bnn_N_Mux_2_2_3_4_4057
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_4_4057_out1 = bnn_Minus_2S_2S_4_960_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4057_out1 = bnn_N_Mux_2_2_3_4_4054_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_4
         always @(s_reg_944 or bnn_Minus_2S_2S_4_960_out1 or bnn_N_Mux_2_2_3_4_4054_in3)
          begin :bnn_N_Mux_2_2_3_4_4060
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_4_4060_out1 = bnn_Minus_2S_2S_4_960_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_4_4060_out1 = bnn_N_Mux_2_2_3_4_4054_in3;
            end
         end

         // resource: mux_2bx2i
         always @(s_reg_959 or bnn_N_Mux_2_2_3_1_3365_out1 or gs_ctrl197)
          begin :drive_bnn_N_Mux_2_2_3_1_4076_in3
            if (gs_ctrl197) begin
               bnn_N_Mux_2_2_3_1_4076_in3 = bnn_N_Mux_2_2_3_1_3365_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4076_in3 = s_reg_959;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_957 or bnn_Minus_2S_2S_1_999_out1 or bnn_N_Mux_2_2_3_1_4076_in3)
          begin :bnn_N_Mux_2_2_3_1_4076
            if (s_reg_957) begin
               bnn_N_Mux_2_2_3_1_4076_out1 = bnn_Minus_2S_2S_1_999_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4076_out1 = bnn_N_Mux_2_2_3_1_4076_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_951 or bnn_Minus_2S_2S_1_999_out1 or bnn_N_Mux_2_2_3_1_4076_in3)
          begin :bnn_N_Mux_2_2_3_1_4078
            if (s_reg_951) begin
               bnn_N_Mux_2_2_3_1_4078_out1 = bnn_Minus_2S_2S_1_999_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4078_out1 = bnn_N_Mux_2_2_3_1_4076_in3;
            end
         end

         // resource: bnn_N_Mux_2_2_3_1
         always @(s_reg_944 or bnn_Minus_2S_2S_1_999_out1 or bnn_N_Mux_2_2_3_1_4076_in3)
          begin :bnn_N_Mux_2_2_3_1_4080
            if (s_reg_944) begin
               bnn_N_Mux_2_2_3_1_4080_out1 = bnn_Minus_2S_2S_1_999_out1;
            end
            else begin
               bnn_N_Mux_2_2_3_1_4080_out1 = bnn_N_Mux_2_2_3_1_4076_in3;
            end
         end

         // resource: bnn_N_Mux_4_2_11_4
         always @(s_reg_1014 or s_reg_1018_slice)
          begin :bnn_N_Mux_4_2_11_4_4090
            if (s_reg_1014) begin
               bnn_N_Mux_4_2_11_4_4090_out1 = {s_reg_1018_slice, 2'd3};
            end
            else begin
               bnn_N_Mux_4_2_11_4_4090_out1 = 4'd00;
            end
         end

         // resource: bnn_N_Mux_4_2_11_4
         always @(s_reg_1015 or s_reg_1018_slice)
          begin :bnn_N_Mux_4_2_11_4_4098
            if (s_reg_1015) begin
               bnn_N_Mux_4_2_11_4_4098_out1 = {s_reg_1018_slice, 2'd3};
            end
            else begin
               bnn_N_Mux_4_2_11_4_4098_out1 = 4'd00;
            end
         end

         // resource: bnn_N_Mux_4_2_11_4
         always @(s_reg_1016 or s_reg_1018_slice)
          begin :bnn_N_Mux_4_2_11_4_4099
            if (s_reg_1016) begin
               bnn_N_Mux_4_2_11_4_4099_out1 = {s_reg_1018_slice, 2'd3};
            end
            else begin
               bnn_N_Mux_4_2_11_4_4099_out1 = 4'd00;
            end
         end

         // resource: bnn_N_Mux_4_2_11_4
         always @(s_reg_870 or s_reg_1018_slice)
          begin :bnn_N_Mux_4_2_11_4_4100
            if (s_reg_870) begin
               bnn_N_Mux_4_2_11_4_4100_out1 = {s_reg_1018_slice, 2'd3};
            end
            else begin
               bnn_N_Mux_4_2_11_4_4100_out1 = 4'd00;
            end
         end

         // resource: bnn_LessThan_10Ux32U_1U_4  instance: bnn_LessThan_10Ux32U_1U_4_4104
         assign bnn_LessThan_10Ux32U_1U_4_4104_out1 = {22'b0000000000000000000000, s_reg_1163} < s_reg_1001;

         // resource: bnn_N_Mux_3_2_6_4
         always @(s_reg_1022 or s_reg_1023)
          begin :bnn_N_Mux_3_2_6_4_4105
            if (s_reg_1023) begin
               bnn_N_Mux_3_2_6_4_4105_out1 = s_reg_1022;
            end
            else begin
               bnn_N_Mux_3_2_6_4_4105_out1 = 3'd0;
            end
         end

         // resource: bnn_Add_2Ux2U_3U_4  instance: bnn_Add_2Ux2U_3U_4_4427
         assign bnn_Add_2Ux2U_3U_4_4427_out1 = {1'b0, s_reg_1004} + 3'd3;

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4430
         assign bnn_Mul_16Sx12S_19S_4_4430_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_1_if_1_dout_wire[11]}}, fixed_buffer_1_if_1_dout_wire};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4433
         assign bnn_Mul_16Sx12S_19S_4_4433_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_2_if_1_dout_wire[11]}}, fixed_buffer_2_if_1_dout_wire};

         // resource: bnn_OrReduction_32U_1U_4  instance: bnn_OrReduction_32U_1U_4_4434
         assign bnn_OrReduction_32U_1U_4_4434_out1 = |s_reg_1002;

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4436
         assign bnn_Mul_16Sx12S_19S_4_4436_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_3_if_1_dout_wire[11]}}, fixed_buffer_3_if_1_dout_wire};

         assign bnn_RightShift_10Ux3U_10U_4_4437_in2 = {s_reg_871[3:0], 6'd00};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4437
         assign bnn_RightShift_10Ux3U_10U_4_4437_out1 = bnn_RightShift_10Ux3U_10U_4_4437_in2 >> {3'b000, s_reg_1012};

         assign bnn_RightShift_10Ux3U_10U_4_4438_in2 = {s_reg_871[3:0], 6'd01};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4438
         assign bnn_RightShift_10Ux3U_10U_4_4438_out1 = bnn_RightShift_10Ux3U_10U_4_4438_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4440
         assign bnn_Mul_16Sx12S_19S_4_4440_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_4_if_1_dout_wire[11]}}, fixed_buffer_4_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4441_in2 = bnn_RightShift_10Ux3U_10U_4_4437_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4441
         assign bnn_LeftShift_9Ux3U_7U_4_4441_out1 = bnn_LeftShift_9Ux3U_7U_4_4441_in2[6:0] << s_reg_1012;

         assign bnn_LeftShift_9Ux3U_7U_4_4442_in2 = bnn_RightShift_10Ux3U_10U_4_4438_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4442
         assign bnn_LeftShift_9Ux3U_7U_4_4442_out1 = bnn_LeftShift_9Ux3U_7U_4_4442_in2[6:0] << s_reg_1012;

         // resource: bnn_N_Mux_6_2_12_4
         always @(bnn_OrReduction_32U_1U_4_4434_out1)
          begin :bnn_N_Mux_6_2_12_4_4443
            if (bnn_OrReduction_32U_1U_4_4434_out1) begin
               bnn_N_Mux_6_2_12_4_4443_out1 = 6'd00;
            end
            else begin
               bnn_N_Mux_6_2_12_4_4443_out1 = 6'd63;
            end
         end

         assign bnn_RightShift_10Ux3U_10U_4_4444_in2 = {s_reg_871[3:0], 6'd02};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4444
         assign bnn_RightShift_10Ux3U_10U_4_4444_out1 = bnn_RightShift_10Ux3U_10U_4_4444_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4446
         assign bnn_Mul_16Sx12S_19S_4_4446_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_5_if_1_dout_wire[11]}}, fixed_buffer_5_if_1_dout_wire};

         assign bnn_LeftShift_1Ux6U_64U_4_4447_in1 = bnn_LeftShift_9Ux3U_7U_4_4441_out1[6:1];

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4447
         assign bnn_LeftShift_1Ux6U_64U_4_4447_out1 = 64'd00000000000000000001 << bnn_LeftShift_1Ux6U_64U_4_4447_in1;

         assign bnn_LeftShift_9Ux3U_7U_4_4449_in2 = bnn_RightShift_10Ux3U_10U_4_4444_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4449
         assign bnn_LeftShift_9Ux3U_7U_4_4449_out1 = bnn_LeftShift_9Ux3U_7U_4_4449_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_2Ux32U_7U_4  instance: bnn_Mod_2Ux32U_7U_4_4450
         assign bnn_Mod_2Ux32U_7U_4_4450_out1 = 2'd2 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4451_in2 = {s_reg_871[3:0], 6'd03};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4451
         assign bnn_RightShift_10Ux3U_10U_4_4451_out1 = bnn_RightShift_10Ux3U_10U_4_4451_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4453
         assign bnn_Mul_16Sx12S_19S_4_4453_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_6_if_1_dout_wire[11]}}, fixed_buffer_6_if_1_dout_wire};

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4454
         assign bnn_NotBit_64U_64U_4_4454_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4447_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4455
         assign bnn_LeftShift_1Ux6U_64U_1_4455_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3375_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4457_in2 = bnn_RightShift_10Ux3U_10U_4_4451_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4457
         assign bnn_LeftShift_9Ux3U_7U_4_4457_out1 = bnn_LeftShift_9Ux3U_7U_4_4457_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_2Ux32U_7U_4  instance: bnn_Mod_2Ux32U_7U_4_4458
         assign bnn_Mod_2Ux32U_7U_4_4458_out1 = 2'd3 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4459_in2 = {s_reg_871[3:0], 6'd04};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4459
         assign bnn_RightShift_10Ux3U_10U_4_4459_out1 = bnn_RightShift_10Ux3U_10U_4_4459_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Equal_2Ux2U_1U_4  instance: bnn_Equal_2Ux2U_1U_4_4460
         assign bnn_Equal_2Ux2U_1U_4_4460_out1 = s_reg_871[1:0] == 2'd3;

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4462
         assign bnn_Mul_16Sx12S_19S_4_4462_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_7_if_1_dout_wire[11]}}, fixed_buffer_7_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4463_ctrl1 = bnn_Add_17Sx16S_17S_1_2389_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4454_out1 or bnn_N_Mux_64_2_2_1_4463_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4463
            if (bnn_N_Mux_64_2_2_1_4463_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4463_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4463_out1 = bnn_NotBit_64U_64U_4_4454_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4464
         assign bnn_NotBit_64U_64U_4_4464_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4455_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4465
         assign bnn_LeftShift_1Ux6U_64U_4_4465_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_4_3070_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4467_in2 = bnn_RightShift_10Ux3U_10U_4_4459_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4467
         assign bnn_LeftShift_9Ux3U_7U_4_4467_out1 = bnn_LeftShift_9Ux3U_7U_4_4467_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_3Ux32U_7U_4  instance: bnn_Mod_3Ux32U_7U_4_4468
         assign bnn_Mod_3Ux32U_7U_4_4468_out1 = 3'd4 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4469_in2 = {s_reg_871[3:0], 6'd05};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4469
         assign bnn_RightShift_10Ux3U_10U_4_4469_out1 = bnn_RightShift_10Ux3U_10U_4_4469_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4471
         assign bnn_Mul_16Sx12S_19S_4_4471_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_8_if_1_dout_wire[11]}}, fixed_buffer_8_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4472
         assign bnn_And_64Sx64S_64S_1_4472_out1 = bnn_N_Mux_64_2_2_1_4463_out1 & Boutword_i0_mi87;

         assign bnn_N_Mux_64_2_2_1_4473_ctrl1 = bnn_Add_17Sx16S_17S_1_3162_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4464_out1 or bnn_N_Mux_64_2_2_1_4473_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4473
            if (bnn_N_Mux_64_2_2_1_4473_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4473_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4473_out1 = bnn_NotBit_64U_64U_4_4464_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4474
         assign bnn_NotBit_64U_64U_4_4474_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4465_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4475
         assign bnn_LeftShift_1Ux6U_64U_4_4475_out1 = 64'd00000000000000000001 << bnn_Add_7Sx6U_7S_4_3098_out1[5:0];

         assign bnn_LeftShift_9Ux3U_7U_4_4477_in2 = bnn_RightShift_10Ux3U_10U_4_4469_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4477
         assign bnn_LeftShift_9Ux3U_7U_4_4477_out1 = bnn_LeftShift_9Ux3U_7U_4_4477_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_3Ux32U_7U_4  instance: bnn_Mod_3Ux32U_7U_4_4478
         assign bnn_Mod_3Ux32U_7U_4_4478_out1 = 3'd5 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4479_in2 = {s_reg_871[3:0], 6'd06};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4479
         assign bnn_RightShift_10Ux3U_10U_4_4479_out1 = bnn_RightShift_10Ux3U_10U_4_4479_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4481
         assign bnn_Mul_16Sx12S_19S_4_4481_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_9_if_1_dout_wire[11]}}, fixed_buffer_9_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4482
         assign bnn_And_64Sx64S_64S_1_4482_out1 = bnn_N_Mux_64_2_2_1_4473_out1 & bnn_And_64Sx64S_64S_1_4472_out1;

         assign bnn_N_Mux_64_2_2_1_4483_ctrl1 = bnn_Add_17Sx16S_17S_1_3118_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4474_out1 or bnn_N_Mux_64_2_2_1_4483_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4483
            if (bnn_N_Mux_64_2_2_1_4483_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4483_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4483_out1 = bnn_NotBit_64U_64U_4_4474_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4484
         assign bnn_NotBit_64U_64U_4_4484_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4475_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4485
         assign bnn_LeftShift_1Ux6U_64U_1_4485_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_407_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4487_in2 = bnn_RightShift_10Ux3U_10U_4_4479_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4487
         assign bnn_LeftShift_9Ux3U_7U_4_4487_out1 = bnn_LeftShift_9Ux3U_7U_4_4487_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_3Ux32U_7U_4  instance: bnn_Mod_3Ux32U_7U_4_4488
         assign bnn_Mod_3Ux32U_7U_4_4488_out1 = 3'd6 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4489_in2 = {s_reg_871[3:0], 6'd07};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4489
         assign bnn_RightShift_10Ux3U_10U_4_4489_out1 = bnn_RightShift_10Ux3U_10U_4_4489_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4491
         assign bnn_Mul_16Sx12S_19S_4_4491_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_10_if_1_dout_wire[11]}}, fixed_buffer_10_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4492
         assign bnn_And_64Sx64S_64S_1_4492_out1 = bnn_N_Mux_64_2_2_1_4483_out1 & bnn_And_64Sx64S_64S_1_4482_out1;

         assign bnn_N_Mux_64_2_2_1_4493_ctrl1 = bnn_Add_17Sx16S_17S_1_3314_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4484_out1 or bnn_N_Mux_64_2_2_1_4493_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4493
            if (bnn_N_Mux_64_2_2_1_4493_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4493_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4493_out1 = bnn_NotBit_64U_64U_4_4484_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4494
         assign bnn_NotBit_64U_64U_4_4494_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4485_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4495
         assign bnn_LeftShift_1Ux6U_64U_1_4495_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_314_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4497_in2 = bnn_RightShift_10Ux3U_10U_4_4489_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4497
         assign bnn_LeftShift_9Ux3U_7U_4_4497_out1 = bnn_LeftShift_9Ux3U_7U_4_4497_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_3Ux32U_7U_4  instance: bnn_Mod_3Ux32U_7U_4_4498
         assign bnn_Mod_3Ux32U_7U_4_4498_out1 = 3'd7 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4499_in2 = {s_reg_871[3:0], 6'd08};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4499
         assign bnn_RightShift_10Ux3U_10U_4_4499_out1 = bnn_RightShift_10Ux3U_10U_4_4499_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4501
         assign bnn_Mul_16Sx12S_19S_4_4501_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_11_if_1_dout_wire[11]}}, fixed_buffer_11_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4502
         assign bnn_And_64Sx64S_64S_1_4502_out1 = bnn_N_Mux_64_2_2_1_4493_out1 & bnn_And_64Sx64S_64S_1_4492_out1;

         assign bnn_N_Mux_64_2_2_1_4503_ctrl1 = bnn_Add_17Sx16S_17S_1_3278_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4494_out1 or bnn_N_Mux_64_2_2_1_4503_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4503
            if (bnn_N_Mux_64_2_2_1_4503_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4503_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4503_out1 = bnn_NotBit_64U_64U_4_4494_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4504
         assign bnn_NotBit_64U_64U_4_4504_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4495_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4505
         assign bnn_LeftShift_1Ux6U_64U_1_4505_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_274_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4507_in2 = bnn_RightShift_10Ux3U_10U_4_4499_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4507
         assign bnn_LeftShift_9Ux3U_7U_4_4507_out1 = bnn_LeftShift_9Ux3U_7U_4_4507_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4508
         assign bnn_Mod_4Ux32U_7U_4_4508_out1 = 4'd08 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4509_in2 = {s_reg_871[3:0], 6'd09};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4509
         assign bnn_RightShift_10Ux3U_10U_4_4509_out1 = bnn_RightShift_10Ux3U_10U_4_4509_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4511
         assign bnn_Mul_16Sx12S_19S_4_4511_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_12_if_1_dout_wire[11]}}, fixed_buffer_12_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4512
         assign bnn_And_64Sx64S_64S_1_4512_out1 = bnn_N_Mux_64_2_2_1_4503_out1 & bnn_And_64Sx64S_64S_1_4502_out1;

         assign bnn_N_Mux_64_2_2_1_4513_ctrl1 = bnn_Add_17Sx16S_17S_1_3247_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4504_out1 or bnn_N_Mux_64_2_2_1_4513_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4513
            if (bnn_N_Mux_64_2_2_1_4513_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4513_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4513_out1 = bnn_NotBit_64U_64U_4_4504_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4514
         assign bnn_NotBit_64U_64U_4_4514_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4505_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4515
         assign bnn_LeftShift_1Ux6U_64U_1_4515_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_282_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4517_in2 = bnn_RightShift_10Ux3U_10U_4_4509_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4517
         assign bnn_LeftShift_9Ux3U_7U_4_4517_out1 = bnn_LeftShift_9Ux3U_7U_4_4517_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4518
         assign bnn_Mod_4Ux32U_7U_4_4518_out1 = 4'd09 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4519_in2 = {s_reg_871[3:0], 6'd10};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4519
         assign bnn_RightShift_10Ux3U_10U_4_4519_out1 = bnn_RightShift_10Ux3U_10U_4_4519_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4521
         assign bnn_Mul_16Sx12S_19S_4_4521_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_13_if_1_dout_wire[11]}}, fixed_buffer_13_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4522
         assign bnn_And_64Sx64S_64S_1_4522_out1 = bnn_N_Mux_64_2_2_1_4513_out1 & bnn_And_64Sx64S_64S_1_4512_out1;

         assign bnn_N_Mux_64_2_2_1_4523_ctrl1 = bnn_Add_17Sx16S_17S_1_3262_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4514_out1 or bnn_N_Mux_64_2_2_1_4523_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4523
            if (bnn_N_Mux_64_2_2_1_4523_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4523_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4523_out1 = bnn_NotBit_64U_64U_4_4514_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4524
         assign bnn_NotBit_64U_64U_4_4524_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4515_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4525
         assign bnn_LeftShift_1Ux6U_64U_1_4525_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_298_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4527_in2 = bnn_RightShift_10Ux3U_10U_4_4519_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4527
         assign bnn_LeftShift_9Ux3U_7U_4_4527_out1 = bnn_LeftShift_9Ux3U_7U_4_4527_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4528
         assign bnn_Mod_4Ux32U_7U_4_4528_out1 = 4'd10 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4529_in2 = {s_reg_871[3:0], 6'd11};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4529
         assign bnn_RightShift_10Ux3U_10U_4_4529_out1 = bnn_RightShift_10Ux3U_10U_4_4529_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4531
         assign bnn_Mul_16Sx12S_19S_4_4531_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_14_if_1_dout_wire[11]}}, fixed_buffer_14_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4532
         assign bnn_And_64Sx64S_64S_1_4532_out1 = bnn_N_Mux_64_2_2_1_4523_out1 & bnn_And_64Sx64S_64S_1_4522_out1;

         assign bnn_N_Mux_64_2_2_1_4533_ctrl1 = bnn_Add_17Sx16S_17S_1_3296_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4524_out1 or bnn_N_Mux_64_2_2_1_4533_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4533
            if (bnn_N_Mux_64_2_2_1_4533_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4533_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4533_out1 = bnn_NotBit_64U_64U_4_4524_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4534
         assign bnn_NotBit_64U_64U_4_4534_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4525_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4535
         assign bnn_LeftShift_1Ux6U_64U_1_4535_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_345_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4537_in2 = bnn_RightShift_10Ux3U_10U_4_4529_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4537
         assign bnn_LeftShift_9Ux3U_7U_4_4537_out1 = bnn_LeftShift_9Ux3U_7U_4_4537_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4538
         assign bnn_Mod_4Ux32U_7U_4_4538_out1 = 4'd11 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4539_in2 = {s_reg_871[3:0], 6'd12};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4539
         assign bnn_RightShift_10Ux3U_10U_4_4539_out1 = bnn_RightShift_10Ux3U_10U_4_4539_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4541
         assign bnn_Mul_16Sx12S_19S_4_4541_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_15_if_1_dout_wire[11]}}, fixed_buffer_15_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4542
         assign bnn_And_64Sx64S_64S_1_4542_out1 = bnn_N_Mux_64_2_2_1_4533_out1 & bnn_And_64Sx64S_64S_1_4532_out1;

         assign bnn_N_Mux_64_2_2_1_4543_ctrl1 = bnn_Add_17Sx16S_17S_1_3097_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4534_out1 or bnn_N_Mux_64_2_2_1_4543_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4543
            if (bnn_N_Mux_64_2_2_1_4543_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4543_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4543_out1 = bnn_NotBit_64U_64U_4_4534_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4544
         assign bnn_NotBit_64U_64U_4_4544_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4535_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4545
         assign bnn_LeftShift_1Ux6U_64U_1_4545_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_365_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4547_in2 = bnn_RightShift_10Ux3U_10U_4_4539_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4547
         assign bnn_LeftShift_9Ux3U_7U_4_4547_out1 = bnn_LeftShift_9Ux3U_7U_4_4547_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4548
         assign bnn_Mod_4Ux32U_7U_4_4548_out1 = 4'd12 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4549_in2 = {s_reg_871[3:0], 6'd13};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4549
         assign bnn_RightShift_10Ux3U_10U_4_4549_out1 = bnn_RightShift_10Ux3U_10U_4_4549_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4551
         assign bnn_Mul_16Sx12S_19S_4_4551_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_16_if_1_dout_wire[11]}}, fixed_buffer_16_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4552
         assign bnn_And_64Sx64S_64S_1_4552_out1 = bnn_N_Mux_64_2_2_1_4543_out1 & bnn_And_64Sx64S_64S_1_4542_out1;

         assign bnn_N_Mux_64_2_2_1_4553_ctrl1 = bnn_Add_17Sx16S_17S_1_3137_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4544_out1 or bnn_N_Mux_64_2_2_1_4553_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4553
            if (bnn_N_Mux_64_2_2_1_4553_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4553_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4553_out1 = bnn_NotBit_64U_64U_4_4544_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4554
         assign bnn_NotBit_64U_64U_4_4554_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4545_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4555
         assign bnn_LeftShift_1Ux6U_64U_1_4555_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_409_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4557_in2 = bnn_RightShift_10Ux3U_10U_4_4549_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4557
         assign bnn_LeftShift_9Ux3U_7U_4_4557_out1 = bnn_LeftShift_9Ux3U_7U_4_4557_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4558
         assign bnn_Mod_4Ux32U_7U_4_4558_out1 = 4'd13 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4559_in2 = {s_reg_871[3:0], 6'd14};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4559
         assign bnn_RightShift_10Ux3U_10U_4_4559_out1 = bnn_RightShift_10Ux3U_10U_4_4559_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4561
         assign bnn_Mul_16Sx12S_19S_4_4561_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_17_if_1_dout_wire[11]}}, fixed_buffer_17_if_1_dout_wire};

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_4562
         assign bnn_And_64Sx64S_64S_1_4562_out1 = bnn_N_Mux_64_2_2_1_4553_out1 & bnn_And_64Sx64S_64S_1_4552_out1;

         assign bnn_N_Mux_64_2_2_1_4563_ctrl1 = bnn_Add_17Sx16S_17S_1_3155_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4554_out1 or bnn_N_Mux_64_2_2_1_4563_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4563
            if (bnn_N_Mux_64_2_2_1_4563_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4563_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4563_out1 = bnn_NotBit_64U_64U_4_4554_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4564
         assign bnn_NotBit_64U_64U_4_4564_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4555_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4565
         assign bnn_LeftShift_1Ux6U_64U_1_4565_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_457_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4567_in2 = bnn_RightShift_10Ux3U_10U_4_4559_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4567
         assign bnn_LeftShift_9Ux3U_7U_4_4567_out1 = bnn_LeftShift_9Ux3U_7U_4_4567_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4568
         assign bnn_Mod_4Ux32U_7U_4_4568_out1 = 4'd14 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4569_in2 = {s_reg_871[3:0], 6'd15};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4569
         assign bnn_RightShift_10Ux3U_10U_4_4569_out1 = bnn_RightShift_10Ux3U_10U_4_4569_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4571
         assign bnn_Mul_16Sx12S_19S_4_4571_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_18_if_1_dout_wire[11]}}, fixed_buffer_18_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4572_ctrl1 = bnn_Add_17Sx16S_17S_1_3174_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4564_out1 or bnn_N_Mux_64_2_2_1_4572_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4572
            if (bnn_N_Mux_64_2_2_1_4572_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4572_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4572_out1 = bnn_NotBit_64U_64U_4_4564_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4573
         assign bnn_NotBit_64U_64U_4_4573_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4565_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4574
         assign bnn_LeftShift_1Ux6U_64U_1_4574_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_699_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4576_in2 = bnn_RightShift_10Ux3U_10U_4_4569_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4576
         assign bnn_LeftShift_9Ux3U_7U_4_4576_out1 = bnn_LeftShift_9Ux3U_7U_4_4576_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_4Ux32U_7U_4  instance: bnn_Mod_4Ux32U_7U_4_4577
         assign bnn_Mod_4Ux32U_7U_4_4577_out1 = 4'd15 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4578_in2 = {s_reg_871[3:0], 6'd16};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4578
         assign bnn_RightShift_10Ux3U_10U_4_4578_out1 = bnn_RightShift_10Ux3U_10U_4_4578_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4580
         assign bnn_Mul_16Sx12S_19S_4_4580_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_19_if_1_dout_wire[11]}}, fixed_buffer_19_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4581_ctrl1 = bnn_Add_17Sx16S_17S_1_3192_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4573_out1 or bnn_N_Mux_64_2_2_1_4581_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4581
            if (bnn_N_Mux_64_2_2_1_4581_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4581_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4581_out1 = bnn_NotBit_64U_64U_4_4573_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4582
         assign bnn_NotBit_64U_64U_4_4582_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4574_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4583
         assign bnn_LeftShift_1Ux6U_64U_1_4583_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_887_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4585_in2 = bnn_RightShift_10Ux3U_10U_4_4578_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4585
         assign bnn_LeftShift_9Ux3U_7U_4_4585_out1 = bnn_LeftShift_9Ux3U_7U_4_4585_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4586
         assign bnn_Mod_5Ux32U_7U_1_4586_out1 = 5'd16 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4587_in2 = {s_reg_871[3:0], 6'd17};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4587
         assign bnn_RightShift_10Ux3U_10U_4_4587_out1 = bnn_RightShift_10Ux3U_10U_4_4587_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4589
         assign bnn_Mul_16Sx12S_19S_4_4589_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_20_if_1_dout_wire[11]}}, fixed_buffer_20_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4590_ctrl1 = bnn_Add_17Sx16S_17S_1_3207_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4582_out1 or bnn_N_Mux_64_2_2_1_4590_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4590
            if (bnn_N_Mux_64_2_2_1_4590_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4590_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4590_out1 = bnn_NotBit_64U_64U_4_4582_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4591
         assign bnn_NotBit_64U_64U_4_4591_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4583_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_4592
         assign bnn_LeftShift_1Ux6U_64U_1_4592_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_1526_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4594_in2 = bnn_RightShift_10Ux3U_10U_4_4587_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4594
         assign bnn_LeftShift_9Ux3U_7U_4_4594_out1 = bnn_LeftShift_9Ux3U_7U_4_4594_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4595
         assign bnn_Mod_5Ux32U_7U_1_4595_out1 = 5'd17 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4596_in2 = {s_reg_871[3:0], 6'd18};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4596
         assign bnn_RightShift_10Ux3U_10U_4_4596_out1 = bnn_RightShift_10Ux3U_10U_4_4596_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4598
         assign bnn_Mul_16Sx12S_19S_4_4598_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_21_if_1_dout_wire[11]}}, fixed_buffer_21_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4599_ctrl1 = bnn_Add_17Sx16S_17S_1_3220_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4591_out1 or bnn_N_Mux_64_2_2_1_4599_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4599
            if (bnn_N_Mux_64_2_2_1_4599_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4599_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4599_out1 = bnn_NotBit_64U_64U_4_4591_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4600
         assign bnn_NotBit_64U_64U_4_4600_out1 = ~bnn_LeftShift_1Ux6U_64U_1_4592_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4601
         assign bnn_LeftShift_1Ux6U_64U_4_4601_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2337_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4603_in2 = bnn_RightShift_10Ux3U_10U_4_4596_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4603
         assign bnn_LeftShift_9Ux3U_7U_4_4603_out1 = bnn_LeftShift_9Ux3U_7U_4_4603_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4604
         assign bnn_Mod_5Ux32U_7U_1_4604_out1 = 5'd18 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4605_in2 = {s_reg_871[3:0], 6'd19};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4605
         assign bnn_RightShift_10Ux3U_10U_4_4605_out1 = bnn_RightShift_10Ux3U_10U_4_4605_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4607
         assign bnn_Mul_16Sx12S_19S_4_4607_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_22_if_1_dout_wire[11]}}, fixed_buffer_22_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4608_ctrl1 = bnn_Add_17Sx16S_17S_1_3233_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4600_out1 or bnn_N_Mux_64_2_2_1_4608_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4608
            if (bnn_N_Mux_64_2_2_1_4608_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4608_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4608_out1 = bnn_NotBit_64U_64U_4_4600_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4609
         assign bnn_NotBit_64U_64U_4_4609_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4601_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4610
         assign bnn_LeftShift_1Ux6U_64U_4_4610_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2362_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4612_in2 = bnn_RightShift_10Ux3U_10U_4_4605_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4612
         assign bnn_LeftShift_9Ux3U_7U_4_4612_out1 = bnn_LeftShift_9Ux3U_7U_4_4612_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4613
         assign bnn_Mod_5Ux32U_7U_1_4613_out1 = 5'd19 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4614_in2 = {s_reg_871[3:0], 6'd20};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4614
         assign bnn_RightShift_10Ux3U_10U_4_4614_out1 = bnn_RightShift_10Ux3U_10U_4_4614_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4616
         assign bnn_Mul_16Sx12S_19S_4_4616_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_23_if_1_dout_wire[11]}}, fixed_buffer_23_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4617_ctrl1 = bnn_Add_17Sx16S_17S_1_3329_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4609_out1 or bnn_N_Mux_64_2_2_1_4617_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4617
            if (bnn_N_Mux_64_2_2_1_4617_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4617_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4617_out1 = bnn_NotBit_64U_64U_4_4609_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4618
         assign bnn_NotBit_64U_64U_4_4618_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4610_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4619
         assign bnn_LeftShift_1Ux6U_64U_4_4619_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2365_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4621_in2 = bnn_RightShift_10Ux3U_10U_4_4614_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4621
         assign bnn_LeftShift_9Ux3U_7U_4_4621_out1 = bnn_LeftShift_9Ux3U_7U_4_4621_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4622
         assign bnn_Mod_5Ux32U_7U_1_4622_out1 = 5'd20 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4623_in2 = {s_reg_871[3:0], 6'd21};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4623
         assign bnn_RightShift_10Ux3U_10U_4_4623_out1 = bnn_RightShift_10Ux3U_10U_4_4623_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4625
         assign bnn_Mul_16Sx12S_19S_4_4625_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_24_if_1_dout_wire[11]}}, fixed_buffer_24_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4626_ctrl1 = bnn_Add_17Sx16S_17S_1_3342_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4618_out1 or bnn_N_Mux_64_2_2_1_4626_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4626
            if (bnn_N_Mux_64_2_2_1_4626_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4626_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4626_out1 = bnn_NotBit_64U_64U_4_4618_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4627
         assign bnn_NotBit_64U_64U_4_4627_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4619_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4628
         assign bnn_LeftShift_1Ux6U_64U_4_4628_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2393_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4630_in2 = bnn_RightShift_10Ux3U_10U_4_4623_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4630
         assign bnn_LeftShift_9Ux3U_7U_4_4630_out1 = bnn_LeftShift_9Ux3U_7U_4_4630_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4631
         assign bnn_Mod_5Ux32U_7U_1_4631_out1 = 5'd21 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4632_in2 = {s_reg_871[3:0], 6'd22};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4632
         assign bnn_RightShift_10Ux3U_10U_4_4632_out1 = bnn_RightShift_10Ux3U_10U_4_4632_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4634
         assign bnn_Mul_16Sx12S_19S_4_4634_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_25_if_1_dout_wire[11]}}, fixed_buffer_25_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4635_ctrl1 = bnn_Add_17Sx16S_17S_1_3355_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4627_out1 or bnn_N_Mux_64_2_2_1_4635_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4635
            if (bnn_N_Mux_64_2_2_1_4635_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4635_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4635_out1 = bnn_NotBit_64U_64U_4_4627_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4636
         assign bnn_NotBit_64U_64U_4_4636_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4628_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4637
         assign bnn_LeftShift_1Ux6U_64U_4_4637_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2420_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4639_in2 = bnn_RightShift_10Ux3U_10U_4_4632_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4639
         assign bnn_LeftShift_9Ux3U_7U_4_4639_out1 = bnn_LeftShift_9Ux3U_7U_4_4639_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4640
         assign bnn_Mod_5Ux32U_7U_1_4640_out1 = 5'd22 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4641_in2 = {s_reg_871[3:0], 6'd23};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4641
         assign bnn_RightShift_10Ux3U_10U_4_4641_out1 = bnn_RightShift_10Ux3U_10U_4_4641_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4643
         assign bnn_Mul_16Sx12S_19S_4_4643_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_26_if_1_dout_wire[11]}}, fixed_buffer_26_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4644_ctrl1 = bnn_Add_17Sx16S_17S_1_3369_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4636_out1 or bnn_N_Mux_64_2_2_1_4644_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4644
            if (bnn_N_Mux_64_2_2_1_4644_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4644_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4644_out1 = bnn_NotBit_64U_64U_4_4636_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4645
         assign bnn_NotBit_64U_64U_4_4645_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4637_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4646
         assign bnn_LeftShift_1Ux6U_64U_4_4646_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2447_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4648_in2 = bnn_RightShift_10Ux3U_10U_4_4641_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4648
         assign bnn_LeftShift_9Ux3U_7U_4_4648_out1 = bnn_LeftShift_9Ux3U_7U_4_4648_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4649
         assign bnn_Mod_5Ux32U_7U_1_4649_out1 = 5'd23 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4650_in2 = {s_reg_871[3:0], 6'd24};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4650
         assign bnn_RightShift_10Ux3U_10U_4_4650_out1 = bnn_RightShift_10Ux3U_10U_4_4650_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4652
         assign bnn_Mul_16Sx12S_19S_4_4652_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_27_if_1_dout_wire[11]}}, fixed_buffer_27_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4653_ctrl1 = bnn_Add_17Sx16S_17S_1_3384_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4645_out1 or bnn_N_Mux_64_2_2_1_4653_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4653
            if (bnn_N_Mux_64_2_2_1_4653_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4653_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4653_out1 = bnn_NotBit_64U_64U_4_4645_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4654
         assign bnn_NotBit_64U_64U_4_4654_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4646_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4655
         assign bnn_LeftShift_1Ux6U_64U_4_4655_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2474_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4657_in2 = bnn_RightShift_10Ux3U_10U_4_4650_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4657
         assign bnn_LeftShift_9Ux3U_7U_4_4657_out1 = bnn_LeftShift_9Ux3U_7U_4_4657_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4658
         assign bnn_Mod_5Ux32U_7U_1_4658_out1 = 5'd24 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4659_in2 = {s_reg_871[3:0], 6'd25};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4659
         assign bnn_RightShift_10Ux3U_10U_4_4659_out1 = bnn_RightShift_10Ux3U_10U_4_4659_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4661
         assign bnn_Mul_16Sx12S_19S_4_4661_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_28_if_1_dout_wire[11]}}, fixed_buffer_28_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4662_ctrl1 = bnn_Add_17Sx16S_17S_1_3400_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4654_out1 or bnn_N_Mux_64_2_2_1_4662_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4662
            if (bnn_N_Mux_64_2_2_1_4662_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4662_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4662_out1 = bnn_NotBit_64U_64U_4_4654_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4663
         assign bnn_NotBit_64U_64U_4_4663_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4655_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4664
         assign bnn_LeftShift_1Ux6U_64U_4_4664_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2501_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4666_in2 = bnn_RightShift_10Ux3U_10U_4_4659_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4666
         assign bnn_LeftShift_9Ux3U_7U_4_4666_out1 = bnn_LeftShift_9Ux3U_7U_4_4666_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4667
         assign bnn_Mod_5Ux32U_7U_1_4667_out1 = 5'd25 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4668_in2 = {s_reg_871[3:0], 6'd26};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4668
         assign bnn_RightShift_10Ux3U_10U_4_4668_out1 = bnn_RightShift_10Ux3U_10U_4_4668_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4670
         assign bnn_Mul_16Sx12S_19S_4_4670_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_29_if_1_dout_wire[11]}}, fixed_buffer_29_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4671_ctrl1 = bnn_Add_17Sx16S_17S_1_3418_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4663_out1 or bnn_N_Mux_64_2_2_1_4671_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4671
            if (bnn_N_Mux_64_2_2_1_4671_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4671_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4671_out1 = bnn_NotBit_64U_64U_4_4663_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4672
         assign bnn_NotBit_64U_64U_4_4672_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4664_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4673
         assign bnn_LeftShift_1Ux6U_64U_4_4673_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2555_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4675_in2 = bnn_RightShift_10Ux3U_10U_4_4668_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4675
         assign bnn_LeftShift_9Ux3U_7U_4_4675_out1 = bnn_LeftShift_9Ux3U_7U_4_4675_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4676
         assign bnn_Mod_5Ux32U_7U_1_4676_out1 = 5'd26 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4677_in2 = {s_reg_871[3:0], 6'd27};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4677
         assign bnn_RightShift_10Ux3U_10U_4_4677_out1 = bnn_RightShift_10Ux3U_10U_4_4677_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4679
         assign bnn_Mul_16Sx12S_19S_4_4679_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_30_if_1_dout_wire[11]}}, fixed_buffer_30_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4680_ctrl1 = bnn_Add_17Sx16S_17S_1_3436_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4672_out1 or bnn_N_Mux_64_2_2_1_4680_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4680
            if (bnn_N_Mux_64_2_2_1_4680_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4680_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4680_out1 = bnn_NotBit_64U_64U_4_4672_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4681
         assign bnn_NotBit_64U_64U_4_4681_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4673_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4682
         assign bnn_LeftShift_1Ux6U_64U_4_4682_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2582_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4684_in2 = bnn_RightShift_10Ux3U_10U_4_4677_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4684
         assign bnn_LeftShift_9Ux3U_7U_4_4684_out1 = bnn_LeftShift_9Ux3U_7U_4_4684_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4685
         assign bnn_Mod_5Ux32U_7U_1_4685_out1 = 5'd27 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4686_in2 = {s_reg_871[3:0], 6'd28};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4686
         assign bnn_RightShift_10Ux3U_10U_4_4686_out1 = bnn_RightShift_10Ux3U_10U_4_4686_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4688
         assign bnn_Mul_16Sx12S_19S_4_4688_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_31_if_1_dout_wire[11]}}, fixed_buffer_31_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4689_ctrl1 = bnn_Add_17Sx16S_17S_1_3451_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4681_out1 or bnn_N_Mux_64_2_2_1_4689_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4689
            if (bnn_N_Mux_64_2_2_1_4689_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4689_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4689_out1 = bnn_NotBit_64U_64U_4_4681_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4690
         assign bnn_NotBit_64U_64U_4_4690_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4682_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4691
         assign bnn_LeftShift_1Ux6U_64U_4_4691_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2609_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4693_in2 = bnn_RightShift_10Ux3U_10U_4_4686_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4693
         assign bnn_LeftShift_9Ux3U_7U_4_4693_out1 = bnn_LeftShift_9Ux3U_7U_4_4693_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4694
         assign bnn_Mod_5Ux32U_7U_1_4694_out1 = 5'd28 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4695_in2 = {s_reg_871[3:0], 6'd29};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4695
         assign bnn_RightShift_10Ux3U_10U_4_4695_out1 = bnn_RightShift_10Ux3U_10U_4_4695_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4697
         assign bnn_Mul_16Sx12S_19S_4_4697_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_32_if_1_dout_wire[11]}}, fixed_buffer_32_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4698_ctrl1 = bnn_Add_17Sx16S_17S_1_3464_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4690_out1 or bnn_N_Mux_64_2_2_1_4698_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4698
            if (bnn_N_Mux_64_2_2_1_4698_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4698_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4698_out1 = bnn_NotBit_64U_64U_4_4690_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4699
         assign bnn_NotBit_64U_64U_4_4699_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4691_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4700
         assign bnn_LeftShift_1Ux6U_64U_4_4700_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2636_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4702_in2 = bnn_RightShift_10Ux3U_10U_4_4695_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4702
         assign bnn_LeftShift_9Ux3U_7U_4_4702_out1 = bnn_LeftShift_9Ux3U_7U_4_4702_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4703
         assign bnn_Mod_5Ux32U_7U_1_4703_out1 = 5'd29 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4704_in2 = {s_reg_871[3:0], 6'd30};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4704
         assign bnn_RightShift_10Ux3U_10U_4_4704_out1 = bnn_RightShift_10Ux3U_10U_4_4704_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4706
         assign bnn_Mul_16Sx12S_19S_4_4706_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_33_if_1_dout_wire[11]}}, fixed_buffer_33_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4707_ctrl1 = bnn_Add_17Sx16S_17S_1_3477_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4699_out1 or bnn_N_Mux_64_2_2_1_4707_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4707
            if (bnn_N_Mux_64_2_2_1_4707_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4707_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4707_out1 = bnn_NotBit_64U_64U_4_4699_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4708
         assign bnn_NotBit_64U_64U_4_4708_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4700_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4709
         assign bnn_LeftShift_1Ux6U_64U_4_4709_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2663_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4711_in2 = bnn_RightShift_10Ux3U_10U_4_4704_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4711
         assign bnn_LeftShift_9Ux3U_7U_4_4711_out1 = bnn_LeftShift_9Ux3U_7U_4_4711_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4712
         assign bnn_Mod_5Ux32U_7U_1_4712_out1 = 5'd30 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4713_in2 = {s_reg_871[3:0], 6'd31};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4713
         assign bnn_RightShift_10Ux3U_10U_4_4713_out1 = bnn_RightShift_10Ux3U_10U_4_4713_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4715
         assign bnn_Mul_16Sx12S_19S_4_4715_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_34_if_1_dout_wire[11]}}, fixed_buffer_34_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4716_ctrl1 = bnn_Add_17Sx16S_17S_1_3491_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4708_out1 or bnn_N_Mux_64_2_2_1_4716_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4716
            if (bnn_N_Mux_64_2_2_1_4716_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4716_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4716_out1 = bnn_NotBit_64U_64U_4_4708_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4717
         assign bnn_NotBit_64U_64U_4_4717_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4709_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4718
         assign bnn_LeftShift_1Ux6U_64U_4_4718_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2690_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4720_in2 = bnn_RightShift_10Ux3U_10U_4_4713_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4720
         assign bnn_LeftShift_9Ux3U_7U_4_4720_out1 = bnn_LeftShift_9Ux3U_7U_4_4720_in2[6:0] << s_reg_1012;

         // resource: bnn_Mod_5Ux32U_7U_1  instance: bnn_Mod_5Ux32U_7U_1_4721
         assign bnn_Mod_5Ux32U_7U_1_4721_out1 = 5'd31 % s_reg_1002;

         assign bnn_RightShift_10Ux3U_10U_4_4722_in2 = {s_reg_871[3:0], 6'd32};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4722
         assign bnn_RightShift_10Ux3U_10U_4_4722_out1 = bnn_RightShift_10Ux3U_10U_4_4722_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4724
         assign bnn_Mul_16Sx12S_19S_4_4724_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_35_if_1_dout_wire[11]}}, fixed_buffer_35_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4725_ctrl1 = bnn_Add_17Sx16S_17S_1_3506_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4717_out1 or bnn_N_Mux_64_2_2_1_4725_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4725
            if (bnn_N_Mux_64_2_2_1_4725_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4725_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4725_out1 = bnn_NotBit_64U_64U_4_4717_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4726
         assign bnn_NotBit_64U_64U_4_4726_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4718_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4727
         assign bnn_LeftShift_1Ux6U_64U_4_4727_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2717_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4729_in2 = bnn_RightShift_10Ux3U_10U_4_4722_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4729
         assign bnn_LeftShift_9Ux3U_7U_4_4729_out1 = bnn_LeftShift_9Ux3U_7U_4_4729_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4730_in2 = {s_reg_871[3:0], 6'd33};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4730
         assign bnn_RightShift_10Ux3U_10U_4_4730_out1 = bnn_RightShift_10Ux3U_10U_4_4730_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4732
         assign bnn_Mul_16Sx12S_19S_4_4732_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_36_if_1_dout_wire[11]}}, fixed_buffer_36_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4733_ctrl1 = bnn_Add_17Sx16S_17S_1_3521_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4726_out1 or bnn_N_Mux_64_2_2_1_4733_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4733
            if (bnn_N_Mux_64_2_2_1_4733_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4733_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4733_out1 = bnn_NotBit_64U_64U_4_4726_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4734
         assign bnn_NotBit_64U_64U_4_4734_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4727_out1;

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_4735
         assign bnn_LeftShift_1Ux6U_64U_4_4735_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2772_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4736_in2 = bnn_RightShift_10Ux3U_10U_4_4730_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4736
         assign bnn_LeftShift_9Ux3U_7U_4_4736_out1 = bnn_LeftShift_9Ux3U_7U_4_4736_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4737_in2 = {s_reg_871[3:0], 6'd34};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4737
         assign bnn_RightShift_10Ux3U_10U_4_4737_out1 = bnn_RightShift_10Ux3U_10U_4_4737_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4739
         assign bnn_Mul_16Sx12S_19S_4_4739_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_37_if_1_dout_wire[11]}}, fixed_buffer_37_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4740_ctrl1 = bnn_Add_17Sx16S_17S_1_3534_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4734_out1 or bnn_N_Mux_64_2_2_1_4740_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4740
            if (bnn_N_Mux_64_2_2_1_4740_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4740_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4740_out1 = bnn_NotBit_64U_64U_4_4734_out1;
            end
         end

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_4741
         assign bnn_NotBit_64U_64U_4_4741_out1 = ~bnn_LeftShift_1Ux6U_64U_4_4735_out1;

         assign bnn_LeftShift_9Ux3U_7U_4_4742_in2 = bnn_RightShift_10Ux3U_10U_4_4737_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4742
         assign bnn_LeftShift_9Ux3U_7U_4_4742_out1 = bnn_LeftShift_9Ux3U_7U_4_4742_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4743_in2 = {s_reg_871[3:0], 6'd35};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4743
         assign bnn_RightShift_10Ux3U_10U_4_4743_out1 = bnn_RightShift_10Ux3U_10U_4_4743_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4745
         assign bnn_Mul_16Sx12S_19S_4_4745_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_38_if_1_dout_wire[11]}}, fixed_buffer_38_if_1_dout_wire};

         assign bnn_N_Mux_64_2_2_1_4746_ctrl1 = bnn_Add_17Sx16S_17S_1_3542_out1[16];

         // resource: bnn_N_Mux_64_2_2_1
         always @(bnn_NotBit_64U_64U_4_4741_out1 or bnn_N_Mux_64_2_2_1_4746_ctrl1)
          begin :bnn_N_Mux_64_2_2_1_4746
            if (bnn_N_Mux_64_2_2_1_4746_ctrl1) begin
               bnn_N_Mux_64_2_2_1_4746_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_4746_out1 = bnn_NotBit_64U_64U_4_4741_out1;
            end
         end

         assign bnn_LeftShift_9Ux3U_7U_4_4747_in2 = bnn_RightShift_10Ux3U_10U_4_4743_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4747
         assign bnn_LeftShift_9Ux3U_7U_4_4747_out1 = bnn_LeftShift_9Ux3U_7U_4_4747_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4748_in2 = {s_reg_871[3:0], 6'd36};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4748
         assign bnn_RightShift_10Ux3U_10U_4_4748_out1 = bnn_RightShift_10Ux3U_10U_4_4748_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4750
         assign bnn_Mul_16Sx12S_19S_4_4750_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_39_if_1_dout_wire[11]}}, fixed_buffer_39_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4751_in2 = bnn_RightShift_10Ux3U_10U_4_4748_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4751
         assign bnn_LeftShift_9Ux3U_7U_4_4751_out1 = bnn_LeftShift_9Ux3U_7U_4_4751_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4752_in2 = {s_reg_871[3:0], 6'd37};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4752
         assign bnn_RightShift_10Ux3U_10U_4_4752_out1 = bnn_RightShift_10Ux3U_10U_4_4752_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4754
         assign bnn_Mul_16Sx12S_19S_4_4754_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_40_if_1_dout_wire[11]}}, fixed_buffer_40_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4755_in2 = bnn_RightShift_10Ux3U_10U_4_4752_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4755
         assign bnn_LeftShift_9Ux3U_7U_4_4755_out1 = bnn_LeftShift_9Ux3U_7U_4_4755_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4756_in2 = {s_reg_871[3:0], 6'd38};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4756
         assign bnn_RightShift_10Ux3U_10U_4_4756_out1 = bnn_RightShift_10Ux3U_10U_4_4756_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4758
         assign bnn_Mul_16Sx12S_19S_4_4758_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_41_if_1_dout_wire[11]}}, fixed_buffer_41_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4759_in2 = bnn_RightShift_10Ux3U_10U_4_4756_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4759
         assign bnn_LeftShift_9Ux3U_7U_4_4759_out1 = bnn_LeftShift_9Ux3U_7U_4_4759_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4760_in2 = {s_reg_871[3:0], 6'd39};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4760
         assign bnn_RightShift_10Ux3U_10U_4_4760_out1 = bnn_RightShift_10Ux3U_10U_4_4760_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4762
         assign bnn_Mul_16Sx12S_19S_4_4762_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_42_if_1_dout_wire[11]}}, fixed_buffer_42_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4763_in2 = bnn_RightShift_10Ux3U_10U_4_4760_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4763
         assign bnn_LeftShift_9Ux3U_7U_4_4763_out1 = bnn_LeftShift_9Ux3U_7U_4_4763_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4764_in2 = {s_reg_871[3:0], 6'd40};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4764
         assign bnn_RightShift_10Ux3U_10U_4_4764_out1 = bnn_RightShift_10Ux3U_10U_4_4764_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4766
         assign bnn_Mul_16Sx12S_19S_4_4766_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_43_if_1_dout_wire[11]}}, fixed_buffer_43_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4767_in2 = bnn_RightShift_10Ux3U_10U_4_4764_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4767
         assign bnn_LeftShift_9Ux3U_7U_4_4767_out1 = bnn_LeftShift_9Ux3U_7U_4_4767_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4768_in2 = {s_reg_871[3:0], 6'd41};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4768
         assign bnn_RightShift_10Ux3U_10U_4_4768_out1 = bnn_RightShift_10Ux3U_10U_4_4768_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4770
         assign bnn_Mul_16Sx12S_19S_4_4770_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_44_if_1_dout_wire[11]}}, fixed_buffer_44_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4771_in2 = bnn_RightShift_10Ux3U_10U_4_4768_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4771
         assign bnn_LeftShift_9Ux3U_7U_4_4771_out1 = bnn_LeftShift_9Ux3U_7U_4_4771_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4772_in2 = {s_reg_871[3:0], 6'd42};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4772
         assign bnn_RightShift_10Ux3U_10U_4_4772_out1 = bnn_RightShift_10Ux3U_10U_4_4772_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4774
         assign bnn_Mul_16Sx12S_19S_4_4774_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_45_if_1_dout_wire[11]}}, fixed_buffer_45_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4775_in2 = bnn_RightShift_10Ux3U_10U_4_4772_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4775
         assign bnn_LeftShift_9Ux3U_7U_4_4775_out1 = bnn_LeftShift_9Ux3U_7U_4_4775_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4776_in2 = {s_reg_871[3:0], 6'd43};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4776
         assign bnn_RightShift_10Ux3U_10U_4_4776_out1 = bnn_RightShift_10Ux3U_10U_4_4776_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4778
         assign bnn_Mul_16Sx12S_19S_4_4778_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_46_if_1_dout_wire[11]}}, fixed_buffer_46_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4779_in2 = bnn_RightShift_10Ux3U_10U_4_4776_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4779
         assign bnn_LeftShift_9Ux3U_7U_4_4779_out1 = bnn_LeftShift_9Ux3U_7U_4_4779_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4780_in2 = {s_reg_871[3:0], 6'd44};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4780
         assign bnn_RightShift_10Ux3U_10U_4_4780_out1 = bnn_RightShift_10Ux3U_10U_4_4780_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4782
         assign bnn_Mul_16Sx12S_19S_4_4782_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_47_if_1_dout_wire[11]}}, fixed_buffer_47_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4783_in2 = bnn_RightShift_10Ux3U_10U_4_4780_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4783
         assign bnn_LeftShift_9Ux3U_7U_4_4783_out1 = bnn_LeftShift_9Ux3U_7U_4_4783_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4784_in2 = {s_reg_871[3:0], 6'd45};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4784
         assign bnn_RightShift_10Ux3U_10U_4_4784_out1 = bnn_RightShift_10Ux3U_10U_4_4784_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4786
         assign bnn_Mul_16Sx12S_19S_4_4786_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_48_if_1_dout_wire[11]}}, fixed_buffer_48_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4787_in2 = bnn_RightShift_10Ux3U_10U_4_4784_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4787
         assign bnn_LeftShift_9Ux3U_7U_4_4787_out1 = bnn_LeftShift_9Ux3U_7U_4_4787_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4788_in2 = {s_reg_871[3:0], 6'd46};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4788
         assign bnn_RightShift_10Ux3U_10U_4_4788_out1 = bnn_RightShift_10Ux3U_10U_4_4788_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4790
         assign bnn_Mul_16Sx12S_19S_4_4790_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_49_if_1_dout_wire[11]}}, fixed_buffer_49_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4791_in2 = bnn_RightShift_10Ux3U_10U_4_4788_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4791
         assign bnn_LeftShift_9Ux3U_7U_4_4791_out1 = bnn_LeftShift_9Ux3U_7U_4_4791_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4792_in2 = {s_reg_871[3:0], 6'd47};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4792
         assign bnn_RightShift_10Ux3U_10U_4_4792_out1 = bnn_RightShift_10Ux3U_10U_4_4792_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4794
         assign bnn_Mul_16Sx12S_19S_4_4794_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_50_if_1_dout_wire[11]}}, fixed_buffer_50_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4795_in2 = bnn_RightShift_10Ux3U_10U_4_4792_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4795
         assign bnn_LeftShift_9Ux3U_7U_4_4795_out1 = bnn_LeftShift_9Ux3U_7U_4_4795_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4796_in2 = {s_reg_871[3:0], 6'd48};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4796
         assign bnn_RightShift_10Ux3U_10U_4_4796_out1 = bnn_RightShift_10Ux3U_10U_4_4796_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4798
         assign bnn_Mul_16Sx12S_19S_4_4798_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_51_if_1_dout_wire[11]}}, fixed_buffer_51_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4799_in2 = bnn_RightShift_10Ux3U_10U_4_4796_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4799
         assign bnn_LeftShift_9Ux3U_7U_4_4799_out1 = bnn_LeftShift_9Ux3U_7U_4_4799_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4800_in2 = {s_reg_871[3:0], 6'd49};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4800
         assign bnn_RightShift_10Ux3U_10U_4_4800_out1 = bnn_RightShift_10Ux3U_10U_4_4800_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4802
         assign bnn_Mul_16Sx12S_19S_4_4802_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_52_if_1_dout_wire[11]}}, fixed_buffer_52_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4803_in2 = bnn_RightShift_10Ux3U_10U_4_4800_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4803
         assign bnn_LeftShift_9Ux3U_7U_4_4803_out1 = bnn_LeftShift_9Ux3U_7U_4_4803_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4804_in2 = {s_reg_871[3:0], 6'd50};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4804
         assign bnn_RightShift_10Ux3U_10U_4_4804_out1 = bnn_RightShift_10Ux3U_10U_4_4804_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4806
         assign bnn_Mul_16Sx12S_19S_4_4806_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_53_if_1_dout_wire[11]}}, fixed_buffer_53_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4807_in2 = bnn_RightShift_10Ux3U_10U_4_4804_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4807
         assign bnn_LeftShift_9Ux3U_7U_4_4807_out1 = bnn_LeftShift_9Ux3U_7U_4_4807_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4808_in2 = {s_reg_871[3:0], 6'd51};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4808
         assign bnn_RightShift_10Ux3U_10U_4_4808_out1 = bnn_RightShift_10Ux3U_10U_4_4808_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4810
         assign bnn_Mul_16Sx12S_19S_4_4810_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_54_if_1_dout_wire[11]}}, fixed_buffer_54_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4811_in2 = bnn_RightShift_10Ux3U_10U_4_4808_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4811
         assign bnn_LeftShift_9Ux3U_7U_4_4811_out1 = bnn_LeftShift_9Ux3U_7U_4_4811_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4812_in2 = {s_reg_871[3:0], 6'd52};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4812
         assign bnn_RightShift_10Ux3U_10U_4_4812_out1 = bnn_RightShift_10Ux3U_10U_4_4812_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4814
         assign bnn_Mul_16Sx12S_19S_4_4814_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_55_if_1_dout_wire[11]}}, fixed_buffer_55_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4815_in2 = bnn_RightShift_10Ux3U_10U_4_4812_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4815
         assign bnn_LeftShift_9Ux3U_7U_4_4815_out1 = bnn_LeftShift_9Ux3U_7U_4_4815_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4816_in2 = {s_reg_871[3:0], 6'd53};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4816
         assign bnn_RightShift_10Ux3U_10U_4_4816_out1 = bnn_RightShift_10Ux3U_10U_4_4816_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4818
         assign bnn_Mul_16Sx12S_19S_4_4818_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_56_if_1_dout_wire[11]}}, fixed_buffer_56_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4819_in2 = bnn_RightShift_10Ux3U_10U_4_4816_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4819
         assign bnn_LeftShift_9Ux3U_7U_4_4819_out1 = bnn_LeftShift_9Ux3U_7U_4_4819_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4820_in2 = {s_reg_871[3:0], 6'd54};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4820
         assign bnn_RightShift_10Ux3U_10U_4_4820_out1 = bnn_RightShift_10Ux3U_10U_4_4820_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4822
         assign bnn_Mul_16Sx12S_19S_4_4822_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_57_if_1_dout_wire[11]}}, fixed_buffer_57_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4823_in2 = bnn_RightShift_10Ux3U_10U_4_4820_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4823
         assign bnn_LeftShift_9Ux3U_7U_4_4823_out1 = bnn_LeftShift_9Ux3U_7U_4_4823_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4824_in2 = {s_reg_871[3:0], 6'd55};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4824
         assign bnn_RightShift_10Ux3U_10U_4_4824_out1 = bnn_RightShift_10Ux3U_10U_4_4824_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4826
         assign bnn_Mul_16Sx12S_19S_4_4826_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_58_if_1_dout_wire[11]}}, fixed_buffer_58_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4827_in2 = bnn_RightShift_10Ux3U_10U_4_4824_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4827
         assign bnn_LeftShift_9Ux3U_7U_4_4827_out1 = bnn_LeftShift_9Ux3U_7U_4_4827_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4828_in2 = {s_reg_871[3:0], 6'd56};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4828
         assign bnn_RightShift_10Ux3U_10U_4_4828_out1 = bnn_RightShift_10Ux3U_10U_4_4828_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4830
         assign bnn_Mul_16Sx12S_19S_4_4830_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_59_if_1_dout_wire[11]}}, fixed_buffer_59_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4831_in2 = bnn_RightShift_10Ux3U_10U_4_4828_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4831
         assign bnn_LeftShift_9Ux3U_7U_4_4831_out1 = bnn_LeftShift_9Ux3U_7U_4_4831_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4832_in2 = {s_reg_871[3:0], 6'd57};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4832
         assign bnn_RightShift_10Ux3U_10U_4_4832_out1 = bnn_RightShift_10Ux3U_10U_4_4832_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4834
         assign bnn_Mul_16Sx12S_19S_4_4834_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_60_if_1_dout_wire[11]}}, fixed_buffer_60_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4835_in2 = bnn_RightShift_10Ux3U_10U_4_4832_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4835
         assign bnn_LeftShift_9Ux3U_7U_4_4835_out1 = bnn_LeftShift_9Ux3U_7U_4_4835_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4836_in2 = {s_reg_871[3:0], 6'd58};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4836
         assign bnn_RightShift_10Ux3U_10U_4_4836_out1 = bnn_RightShift_10Ux3U_10U_4_4836_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4838
         assign bnn_Mul_16Sx12S_19S_4_4838_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_61_if_1_dout_wire[11]}}, fixed_buffer_61_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4839_in2 = bnn_RightShift_10Ux3U_10U_4_4836_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4839
         assign bnn_LeftShift_9Ux3U_7U_4_4839_out1 = bnn_LeftShift_9Ux3U_7U_4_4839_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4840_in2 = {s_reg_871[3:0], 6'd59};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4840
         assign bnn_RightShift_10Ux3U_10U_4_4840_out1 = bnn_RightShift_10Ux3U_10U_4_4840_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4842
         assign bnn_Mul_16Sx12S_19S_4_4842_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_62_if_1_dout_wire[11]}}, fixed_buffer_62_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4843_in2 = bnn_RightShift_10Ux3U_10U_4_4840_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4843
         assign bnn_LeftShift_9Ux3U_7U_4_4843_out1 = bnn_LeftShift_9Ux3U_7U_4_4843_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4844_in2 = {s_reg_871[3:0], 6'd60};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4844
         assign bnn_RightShift_10Ux3U_10U_4_4844_out1 = bnn_RightShift_10Ux3U_10U_4_4844_in2 >> {3'b000, s_reg_1012};

         // resource: bnn_Mul_16Sx12S_19S_4  instance: bnn_Mul_16Sx12S_19S_4_4846
         assign bnn_Mul_16Sx12S_19S_4_4846_out1 = {{ 3 {s_reg_1003[15]}}, s_reg_1003[15:0]}*{{ 7 {fixed_buffer_63_if_1_dout_wire[11]}}, fixed_buffer_63_if_1_dout_wire};

         assign bnn_LeftShift_9Ux3U_7U_4_4847_in2 = bnn_RightShift_10Ux3U_10U_4_4844_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4847
         assign bnn_LeftShift_9Ux3U_7U_4_4847_out1 = bnn_LeftShift_9Ux3U_7U_4_4847_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4848_in2 = {s_reg_871[3:0], 6'd61};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4848
         assign bnn_RightShift_10Ux3U_10U_4_4848_out1 = bnn_RightShift_10Ux3U_10U_4_4848_in2 >> {3'b000, s_reg_1012};

         assign bnn_LeftShift_9Ux3U_7U_4_4850_in2 = bnn_RightShift_10Ux3U_10U_4_4848_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4850
         assign bnn_LeftShift_9Ux3U_7U_4_4850_out1 = bnn_LeftShift_9Ux3U_7U_4_4850_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4851_in2 = {s_reg_871[3:0], 6'd62};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4851
         assign bnn_RightShift_10Ux3U_10U_4_4851_out1 = bnn_RightShift_10Ux3U_10U_4_4851_in2 >> {3'b000, s_reg_1012};

         assign bnn_LeftShift_9Ux3U_7U_4_4852_in2 = bnn_RightShift_10Ux3U_10U_4_4851_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4852
         assign bnn_LeftShift_9Ux3U_7U_4_4852_out1 = bnn_LeftShift_9Ux3U_7U_4_4852_in2[6:0] << s_reg_1012;

         assign bnn_RightShift_10Ux3U_10U_4_4853_in2 = {s_reg_871[3:0], 6'd63};

         // resource: bnn_RightShift_10Ux3U_10U_4  instance: bnn_RightShift_10Ux3U_10U_4_4853
         assign bnn_RightShift_10Ux3U_10U_4_4853_out1 = bnn_RightShift_10Ux3U_10U_4_4853_in2 >> {3'b000, s_reg_1012};

         assign bnn_LeftShift_9Ux3U_7U_4_4854_in2 = bnn_RightShift_10Ux3U_10U_4_4853_out1[9:1];

         // resource: bnn_LeftShift_9Ux3U_7U_4  instance: bnn_LeftShift_9Ux3U_7U_4_4854
         assign bnn_LeftShift_9Ux3U_7U_4_4854_out1 = bnn_LeftShift_9Ux3U_7U_4_4854_in2[6:0] << s_reg_1012;

         assign bnn_Mod_6Ux32U_7U_4_4988_in2 = 6'd63;

         assign bnn_Mod_6Ux32U_7U_4_4989_in2 = 6'd62;

         assign bnn_Mod_6Ux32U_7U_4_4990_in2 = 6'd61;

         assign bnn_Mod_6Ux32U_7U_4_4991_in2 = 6'd60;

         assign bnn_Mod_6Ux32U_7U_4_4992_in2 = 6'd59;

         assign bnn_Mod_6Ux32U_7U_4_4993_in2 = 6'd58;

         assign bnn_Mod_6Ux32U_7U_4_4994_in2 = 6'd57;

         assign bnn_Mod_6Ux32U_7U_4_4995_in2 = 6'd56;

         assign bnn_Mod_6Ux32U_7U_4_4996_in2 = 6'd55;

         assign bnn_Mod_6Ux32U_7U_4_4997_in2 = 6'd54;

         assign bnn_Mod_6Ux32U_7U_4_4998_in2 = 6'd53;

         assign bnn_Mod_6Ux32U_7U_4_4999_in2 = 6'd52;

         assign bnn_Mod_6Ux32U_7U_4_5000_in2 = 6'd51;

         assign bnn_Mod_6Ux32U_7U_4_5001_in2 = 6'd50;

         assign bnn_Mod_6Ux32U_7U_4_5002_in2 = 6'd49;

         assign bnn_Mod_6Ux32U_7U_4_5003_in2 = 6'd48;

         assign bnn_Mod_6Ux32U_7U_4_5004_in2 = 6'd47;

         assign bnn_Mod_6Ux32U_7U_4_5005_in2 = 6'd46;

         assign bnn_Mod_6Ux32U_7U_4_5006_in2 = 6'd45;

         assign bnn_Mod_6Ux32U_7U_4_5007_in2 = 6'd44;

         assign bnn_Mod_6Ux32U_7U_4_5008_in2 = 6'd43;

         assign bnn_Mod_6Ux32U_7U_4_5009_in2 = 6'd42;

         assign bnn_Mod_6Ux32U_7U_4_5010_in2 = 6'd41;

         assign bnn_Mod_6Ux32U_7U_4_5011_in2 = 6'd40;

         assign bnn_Mod_6Ux32U_7U_4_5012_in2 = 6'd39;

         assign bnn_Mod_6Ux32U_7U_4_5013_in2 = 6'd38;

         assign bnn_Mod_6Ux32U_7U_4_5014_in2 = 6'd37;

         assign bnn_Mod_6Ux32U_7U_4_5015_in2 = 6'd36;

         assign bnn_Mod_6Ux32U_7U_4_5016_in2 = 6'd35;

         assign bnn_Mod_6Ux32U_7U_4_5017_in2 = 6'd34;

         assign bnn_Mod_6Ux32U_7U_4_5018_in2 = 6'd33;

         assign bnn_Mod_6Ux32U_7U_4_5019_in2 = 6'd32;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5020
         assign bnn_And_64Sx64S_64S_4_5020_out1 = s_reg_1144 & s_reg_897;

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5022
         assign bnn_LeftShift_1Ux6U_64U_1_5022_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3214_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5023
         assign bnn_NotBit_64U_64U_4_5023_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5022_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1060 or bnn_NotBit_64U_64U_4_5023_out1)
          begin :bnn_N_Mux_64_2_2_1_5024
            if (s_reg_1060) begin
               bnn_N_Mux_64_2_2_1_5024_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5024_out1 = bnn_NotBit_64U_64U_4_5023_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_5026
         assign bnn_LeftShift_1Ux6U_64U_4_5026_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3336_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5027
         assign bnn_NotBit_64U_64U_4_5027_out1 = ~bnn_LeftShift_1Ux6U_64U_4_5026_out1;

         // resource: bnn_N_Mux_64_2_2_4
         always @(s_reg_1059 or bnn_NotBit_64U_64U_4_5027_out1)
          begin :bnn_N_Mux_64_2_2_4_5028
            if (s_reg_1059) begin
               bnn_N_Mux_64_2_2_4_5028_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_4_5028_out1 = bnn_NotBit_64U_64U_4_5027_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5030
         assign bnn_LeftShift_1Ux6U_64U_1_5030_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3458_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5031
         assign bnn_NotBit_64U_64U_4_5031_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5030_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1055 or bnn_NotBit_64U_64U_4_5031_out1)
          begin :bnn_N_Mux_64_2_2_1_5032
            if (s_reg_1055) begin
               bnn_N_Mux_64_2_2_1_5032_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5032_out1 = bnn_NotBit_64U_64U_4_5031_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5034
         assign bnn_LeftShift_1Ux6U_64U_1_5034_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_2312_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5035
         assign bnn_NotBit_64U_64U_4_5035_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5034_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1057 or bnn_NotBit_64U_64U_4_5035_out1)
          begin :bnn_N_Mux_64_2_2_1_5036
            if (s_reg_1057) begin
               bnn_N_Mux_64_2_2_1_5036_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5036_out1 = bnn_NotBit_64U_64U_4_5035_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5038
         assign bnn_LeftShift_1Ux6U_64U_1_5038_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3119_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5039
         assign bnn_NotBit_64U_64U_4_5039_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5038_out1;

         // resource: bnn_N_Mux_64_2_2_4
         always @(s_reg_1056 or bnn_NotBit_64U_64U_4_5039_out1)
          begin :bnn_N_Mux_64_2_2_4_5040
            if (s_reg_1056) begin
               bnn_N_Mux_64_2_2_4_5040_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_4_5040_out1 = bnn_NotBit_64U_64U_4_5039_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5042
         assign bnn_LeftShift_1Ux6U_64U_1_5042_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3138_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5043
         assign bnn_NotBit_64U_64U_4_5043_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5042_out1;

         // resource: bnn_N_Mux_64_2_2_4
         always @(s_reg_1054 or bnn_NotBit_64U_64U_4_5043_out1)
          begin :bnn_N_Mux_64_2_2_4_5044
            if (s_reg_1054) begin
               bnn_N_Mux_64_2_2_4_5044_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_4_5044_out1 = bnn_NotBit_64U_64U_4_5043_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5046
         assign bnn_LeftShift_1Ux6U_64U_1_5046_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3156_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5047
         assign bnn_NotBit_64U_64U_4_5047_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5046_out1;

         // resource: bnn_N_Mux_64_2_2_4
         always @(s_reg_1053 or bnn_NotBit_64U_64U_4_5047_out1)
          begin :bnn_N_Mux_64_2_2_4_5048
            if (s_reg_1053) begin
               bnn_N_Mux_64_2_2_4_5048_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_4_5048_out1 = bnn_NotBit_64U_64U_4_5047_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_5050
         assign bnn_LeftShift_1Ux6U_64U_4_5050_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3175_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5051
         assign bnn_NotBit_64U_64U_4_5051_out1 = ~bnn_LeftShift_1Ux6U_64U_4_5050_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1051 or bnn_NotBit_64U_64U_4_5051_out1)
          begin :bnn_N_Mux_64_2_2_1_5052
            if (s_reg_1051) begin
               bnn_N_Mux_64_2_2_1_5052_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5052_out1 = bnn_NotBit_64U_64U_4_5051_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_5054
         assign bnn_LeftShift_1Ux6U_64U_4_5054_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3193_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5055
         assign bnn_NotBit_64U_64U_4_5055_out1 = ~bnn_LeftShift_1Ux6U_64U_4_5054_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1049 or bnn_NotBit_64U_64U_4_5055_out1)
          begin :bnn_N_Mux_64_2_2_1_5056
            if (s_reg_1049) begin
               bnn_N_Mux_64_2_2_1_5056_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5056_out1 = bnn_NotBit_64U_64U_4_5055_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_4  instance: bnn_LeftShift_1Ux6U_64U_4_5058
         assign bnn_LeftShift_1Ux6U_64U_4_5058_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3197_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5059
         assign bnn_NotBit_64U_64U_4_5059_out1 = ~bnn_LeftShift_1Ux6U_64U_4_5058_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1045 or bnn_NotBit_64U_64U_4_5059_out1)
          begin :bnn_N_Mux_64_2_2_1_5060
            if (s_reg_1045) begin
               bnn_N_Mux_64_2_2_1_5060_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5060_out1 = bnn_NotBit_64U_64U_4_5059_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5062
         assign bnn_LeftShift_1Ux6U_64U_1_5062_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3315_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5063
         assign bnn_NotBit_64U_64U_4_5063_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5062_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1042 or bnn_NotBit_64U_64U_4_5063_out1)
          begin :bnn_N_Mux_64_2_2_1_5064
            if (s_reg_1042) begin
               bnn_N_Mux_64_2_2_1_5064_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5064_out1 = bnn_NotBit_64U_64U_4_5063_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5066
         assign bnn_LeftShift_1Ux6U_64U_1_5066_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3319_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5067
         assign bnn_NotBit_64U_64U_4_5067_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5066_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1040 or bnn_NotBit_64U_64U_4_5067_out1)
          begin :bnn_N_Mux_64_2_2_1_5068
            if (s_reg_1040) begin
               bnn_N_Mux_64_2_2_1_5068_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5068_out1 = bnn_NotBit_64U_64U_4_5067_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5070
         assign bnn_LeftShift_1Ux6U_64U_1_5070_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3356_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5071
         assign bnn_NotBit_64U_64U_4_5071_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5070_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1038 or bnn_NotBit_64U_64U_4_5071_out1)
          begin :bnn_N_Mux_64_2_2_1_5072
            if (s_reg_1038) begin
               bnn_N_Mux_64_2_2_1_5072_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5072_out1 = bnn_NotBit_64U_64U_4_5071_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5074
         assign bnn_LeftShift_1Ux6U_64U_1_5074_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3370_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5075
         assign bnn_NotBit_64U_64U_4_5075_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5074_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1037 or bnn_NotBit_64U_64U_4_5075_out1)
          begin :bnn_N_Mux_64_2_2_1_5076
            if (s_reg_1037) begin
               bnn_N_Mux_64_2_2_1_5076_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5076_out1 = bnn_NotBit_64U_64U_4_5075_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5078
         assign bnn_LeftShift_1Ux6U_64U_1_5078_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3385_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5079
         assign bnn_NotBit_64U_64U_4_5079_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5078_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1052 or bnn_NotBit_64U_64U_4_5079_out1)
          begin :bnn_N_Mux_64_2_2_1_5080
            if (s_reg_1052) begin
               bnn_N_Mux_64_2_2_1_5080_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5080_out1 = bnn_NotBit_64U_64U_4_5079_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5082
         assign bnn_LeftShift_1Ux6U_64U_1_5082_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3401_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5083
         assign bnn_NotBit_64U_64U_4_5083_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5082_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1050 or bnn_NotBit_64U_64U_4_5083_out1)
          begin :bnn_N_Mux_64_2_2_1_5084
            if (s_reg_1050) begin
               bnn_N_Mux_64_2_2_1_5084_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5084_out1 = bnn_NotBit_64U_64U_4_5083_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5086
         assign bnn_LeftShift_1Ux6U_64U_1_5086_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3419_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5087
         assign bnn_NotBit_64U_64U_4_5087_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5086_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1048 or bnn_NotBit_64U_64U_4_5087_out1)
          begin :bnn_N_Mux_64_2_2_1_5088
            if (s_reg_1048) begin
               bnn_N_Mux_64_2_2_1_5088_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5088_out1 = bnn_NotBit_64U_64U_4_5087_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5090
         assign bnn_LeftShift_1Ux6U_64U_1_5090_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3437_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5091
         assign bnn_NotBit_64U_64U_4_5091_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5090_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1044 or bnn_NotBit_64U_64U_4_5091_out1)
          begin :bnn_N_Mux_64_2_2_1_5092
            if (s_reg_1044) begin
               bnn_N_Mux_64_2_2_1_5092_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5092_out1 = bnn_NotBit_64U_64U_4_5091_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5094
         assign bnn_LeftShift_1Ux6U_64U_1_5094_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3441_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5095
         assign bnn_NotBit_64U_64U_4_5095_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5094_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1024 or bnn_NotBit_64U_64U_4_5095_out1)
          begin :bnn_N_Mux_64_2_2_1_5096
            if (s_reg_1024) begin
               bnn_N_Mux_64_2_2_1_5096_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5096_out1 = bnn_NotBit_64U_64U_4_5095_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5098
         assign bnn_LeftShift_1Ux6U_64U_1_5098_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3478_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5099
         assign bnn_NotBit_64U_64U_4_5099_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5098_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1023 or bnn_NotBit_64U_64U_4_5099_out1)
          begin :bnn_N_Mux_64_2_2_1_5100
            if (s_reg_1023) begin
               bnn_N_Mux_64_2_2_1_5100_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5100_out1 = bnn_NotBit_64U_64U_4_5099_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5102
         assign bnn_LeftShift_1Ux6U_64U_1_5102_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3492_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5103
         assign bnn_NotBit_64U_64U_4_5103_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5102_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1016 or bnn_NotBit_64U_64U_4_5103_out1)
          begin :bnn_N_Mux_64_2_2_1_5104
            if (s_reg_1016) begin
               bnn_N_Mux_64_2_2_1_5104_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5104_out1 = bnn_NotBit_64U_64U_4_5103_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5106
         assign bnn_LeftShift_1Ux6U_64U_1_5106_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3507_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5107
         assign bnn_NotBit_64U_64U_4_5107_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5106_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1015 or bnn_NotBit_64U_64U_4_5107_out1)
          begin :bnn_N_Mux_64_2_2_1_5108
            if (s_reg_1015) begin
               bnn_N_Mux_64_2_2_1_5108_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5108_out1 = bnn_NotBit_64U_64U_4_5107_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5110
         assign bnn_LeftShift_1Ux6U_64U_1_5110_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3522_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5111
         assign bnn_NotBit_64U_64U_4_5111_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5110_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_1014 or bnn_NotBit_64U_64U_4_5111_out1)
          begin :bnn_N_Mux_64_2_2_1_5112
            if (s_reg_1014) begin
               bnn_N_Mux_64_2_2_1_5112_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5112_out1 = bnn_NotBit_64U_64U_4_5111_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5114
         assign bnn_LeftShift_1Ux6U_64U_1_5114_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3535_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5115
         assign bnn_NotBit_64U_64U_4_5115_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5114_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_957 or bnn_NotBit_64U_64U_4_5115_out1)
          begin :bnn_N_Mux_64_2_2_1_5116
            if (s_reg_957) begin
               bnn_N_Mux_64_2_2_1_5116_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5116_out1 = bnn_NotBit_64U_64U_4_5115_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5118
         assign bnn_LeftShift_1Ux6U_64U_1_5118_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3543_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5119
         assign bnn_NotBit_64U_64U_4_5119_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5118_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_951 or bnn_NotBit_64U_64U_4_5119_out1)
          begin :bnn_N_Mux_64_2_2_1_5120
            if (s_reg_951) begin
               bnn_N_Mux_64_2_2_1_5120_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5120_out1 = bnn_NotBit_64U_64U_4_5119_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5122
         assign bnn_LeftShift_1Ux6U_64U_1_5122_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3234_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5123
         assign bnn_NotBit_64U_64U_4_5123_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5122_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_944 or bnn_NotBit_64U_64U_4_5123_out1)
          begin :bnn_N_Mux_64_2_2_1_5124
            if (s_reg_944) begin
               bnn_N_Mux_64_2_2_1_5124_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5124_out1 = bnn_NotBit_64U_64U_4_5123_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5126
         assign bnn_LeftShift_1Ux6U_64U_1_5126_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3248_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5127
         assign bnn_NotBit_64U_64U_4_5127_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5126_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_939 or bnn_NotBit_64U_64U_4_5127_out1)
          begin :bnn_N_Mux_64_2_2_1_5128
            if (s_reg_939) begin
               bnn_N_Mux_64_2_2_1_5128_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5128_out1 = bnn_NotBit_64U_64U_4_5127_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5130
         assign bnn_LeftShift_1Ux6U_64U_1_5130_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3263_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5131
         assign bnn_NotBit_64U_64U_4_5131_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5130_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_932 or bnn_NotBit_64U_64U_4_5131_out1)
          begin :bnn_N_Mux_64_2_2_1_5132
            if (s_reg_932) begin
               bnn_N_Mux_64_2_2_1_5132_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5132_out1 = bnn_NotBit_64U_64U_4_5131_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5134
         assign bnn_LeftShift_1Ux6U_64U_1_5134_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3279_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5135
         assign bnn_NotBit_64U_64U_4_5135_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5134_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_924 or bnn_NotBit_64U_64U_4_5135_out1)
          begin :bnn_N_Mux_64_2_2_1_5136
            if (s_reg_924) begin
               bnn_N_Mux_64_2_2_1_5136_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5136_out1 = bnn_NotBit_64U_64U_4_5135_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5138
         assign bnn_LeftShift_1Ux6U_64U_1_5138_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3297_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5139
         assign bnn_NotBit_64U_64U_4_5139_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5138_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_916 or bnn_NotBit_64U_64U_4_5139_out1)
          begin :bnn_N_Mux_64_2_2_1_5140
            if (s_reg_916) begin
               bnn_N_Mux_64_2_2_1_5140_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5140_out1 = bnn_NotBit_64U_64U_4_5139_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5142
         assign bnn_LeftShift_1Ux6U_64U_1_5142_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3544_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5143
         assign bnn_NotBit_64U_64U_4_5143_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5142_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_908 or bnn_NotBit_64U_64U_4_5143_out1)
          begin :bnn_N_Mux_64_2_2_1_5144
            if (s_reg_908) begin
               bnn_N_Mux_64_2_2_1_5144_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5144_out1 = bnn_NotBit_64U_64U_4_5143_out1;
            end
         end

         // resource: bnn_LeftShift_1Ux6U_64U_1  instance: bnn_LeftShift_1Ux6U_64U_1_5146
         assign bnn_LeftShift_1Ux6U_64U_1_5146_out1 = 64'd00000000000000000001 << bnn_Add_6Ux6U_6U_1_3199_out1;

         // resource: bnn_NotBit_64U_64U_4  instance: bnn_NotBit_64U_64U_4_5147
         assign bnn_NotBit_64U_64U_4_5147_out1 = ~bnn_LeftShift_1Ux6U_64U_1_5146_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_870 or bnn_NotBit_64U_64U_4_5147_out1)
          begin :bnn_N_Mux_64_2_2_1_5148
            if (s_reg_870) begin
               bnn_N_Mux_64_2_2_1_5148_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5148_out1 = bnn_NotBit_64U_64U_4_5147_out1;
            end
         end

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5149
         assign bnn_And_64Sx64S_64S_4_5149_out1 = s_reg_1145 & bnn_And_64Sx64S_64S_4_5020_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5150
         assign bnn_And_64Sx64S_64S_4_5150_out1 = s_reg_1146 & bnn_And_64Sx64S_64S_4_5149_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5151
         assign bnn_And_64Sx64S_64S_4_5151_out1 = s_reg_1147 & bnn_And_64Sx64S_64S_4_5150_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5152
         assign bnn_And_64Sx64S_64S_4_5152_out1 = s_reg_1148 & bnn_And_64Sx64S_64S_4_5151_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5153
         assign bnn_And_64Sx64S_64S_4_5153_out1 = s_reg_1149 & bnn_And_64Sx64S_64S_4_5152_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5154
         assign bnn_And_64Sx64S_64S_4_5154_out1 = s_reg_1150 & bnn_And_64Sx64S_64S_4_5153_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5155
         assign bnn_And_64Sx64S_64S_4_5155_out1 = s_reg_1151 & bnn_And_64Sx64S_64S_4_5154_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5156
         assign bnn_And_64Sx64S_64S_4_5156_out1 = s_reg_1152 & bnn_And_64Sx64S_64S_4_5155_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5157
         assign bnn_And_64Sx64S_64S_4_5157_out1 = s_reg_1153 & bnn_And_64Sx64S_64S_4_5156_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5158
         assign bnn_And_64Sx64S_64S_4_5158_out1 = s_reg_1154 & bnn_And_64Sx64S_64S_4_5157_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5159
         assign bnn_And_64Sx64S_64S_4_5159_out1 = s_reg_1155 & bnn_And_64Sx64S_64S_4_5158_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5160
         assign bnn_And_64Sx64S_64S_4_5160_out1 = s_reg_1156 & bnn_And_64Sx64S_64S_4_5159_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5161
         assign bnn_And_64Sx64S_64S_4_5161_out1 = s_reg_1157 & bnn_And_64Sx64S_64S_4_5160_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5162
         assign bnn_And_64Sx64S_64S_4_5162_out1 = s_reg_1158 & bnn_And_64Sx64S_64S_4_5161_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5163
         assign bnn_And_64Sx64S_64S_4_5163_out1 = s_reg_1159 & bnn_And_64Sx64S_64S_4_5162_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5164
         assign bnn_And_64Sx64S_64S_4_5164_out1 = s_reg_1160 & bnn_And_64Sx64S_64S_4_5163_out1;

         // resource: bnn_And_64Sx64S_64S_4  instance: bnn_And_64Sx64S_64S_4_5165
         assign bnn_And_64Sx64S_64S_4_5165_out1 = s_reg_1161 & bnn_And_64Sx64S_64S_4_5164_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5166
         assign bnn_And_64Sx64S_64S_1_5166_out1 = s_reg_1162 & bnn_And_64Sx64S_64S_4_5165_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5167
         assign bnn_And_64Sx64S_64S_1_5167_out1 = s_reg_1164 & bnn_And_64Sx64S_64S_1_5166_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5168
         assign bnn_And_64Sx64S_64S_1_5168_out1 = s_reg_1165 & bnn_And_64Sx64S_64S_1_5167_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5169
         assign bnn_And_64Sx64S_64S_1_5169_out1 = s_reg_1166 & bnn_And_64Sx64S_64S_1_5168_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5170
         assign bnn_And_64Sx64S_64S_1_5170_out1 = bnn_N_Mux_64_2_2_1_5148_out1 & bnn_And_64Sx64S_64S_1_5169_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5171
         assign bnn_And_64Sx64S_64S_1_5171_out1 = bnn_N_Mux_64_2_2_1_5144_out1 & bnn_And_64Sx64S_64S_1_5170_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5172
         assign bnn_And_64Sx64S_64S_1_5172_out1 = bnn_N_Mux_64_2_2_1_5140_out1 & bnn_And_64Sx64S_64S_1_5171_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5173
         assign bnn_And_64Sx64S_64S_1_5173_out1 = bnn_N_Mux_64_2_2_1_5136_out1 & bnn_And_64Sx64S_64S_1_5172_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5174
         assign bnn_And_64Sx64S_64S_1_5174_out1 = bnn_N_Mux_64_2_2_1_5132_out1 & bnn_And_64Sx64S_64S_1_5173_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5175
         assign bnn_And_64Sx64S_64S_1_5175_out1 = bnn_N_Mux_64_2_2_1_5128_out1 & bnn_And_64Sx64S_64S_1_5174_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5176
         assign bnn_And_64Sx64S_64S_1_5176_out1 = bnn_N_Mux_64_2_2_1_5124_out1 & bnn_And_64Sx64S_64S_1_5175_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5177
         assign bnn_And_64Sx64S_64S_1_5177_out1 = bnn_N_Mux_64_2_2_1_5120_out1 & bnn_And_64Sx64S_64S_1_5176_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5178
         assign bnn_And_64Sx64S_64S_1_5178_out1 = bnn_N_Mux_64_2_2_1_5116_out1 & bnn_And_64Sx64S_64S_1_5177_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5179
         assign bnn_And_64Sx64S_64S_1_5179_out1 = bnn_N_Mux_64_2_2_1_5112_out1 & bnn_And_64Sx64S_64S_1_5178_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5180
         assign bnn_And_64Sx64S_64S_1_5180_out1 = bnn_N_Mux_64_2_2_1_5108_out1 & bnn_And_64Sx64S_64S_1_5179_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5181
         assign bnn_And_64Sx64S_64S_1_5181_out1 = bnn_N_Mux_64_2_2_1_5104_out1 & bnn_And_64Sx64S_64S_1_5180_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5182
         assign bnn_And_64Sx64S_64S_1_5182_out1 = bnn_N_Mux_64_2_2_1_5100_out1 & bnn_And_64Sx64S_64S_1_5181_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5183
         assign bnn_And_64Sx64S_64S_1_5183_out1 = bnn_N_Mux_64_2_2_1_5096_out1 & bnn_And_64Sx64S_64S_1_5182_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5184
         assign bnn_And_64Sx64S_64S_1_5184_out1 = bnn_N_Mux_64_2_2_1_5092_out1 & bnn_And_64Sx64S_64S_1_5183_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5185
         assign bnn_And_64Sx64S_64S_1_5185_out1 = bnn_N_Mux_64_2_2_1_5088_out1 & bnn_And_64Sx64S_64S_1_5184_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5186
         assign bnn_And_64Sx64S_64S_1_5186_out1 = bnn_N_Mux_64_2_2_1_5084_out1 & bnn_And_64Sx64S_64S_1_5185_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5187
         assign bnn_And_64Sx64S_64S_1_5187_out1 = bnn_N_Mux_64_2_2_1_5080_out1 & bnn_And_64Sx64S_64S_1_5186_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5188
         assign bnn_And_64Sx64S_64S_1_5188_out1 = bnn_N_Mux_64_2_2_1_5076_out1 & bnn_And_64Sx64S_64S_1_5187_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5189
         assign bnn_And_64Sx64S_64S_1_5189_out1 = bnn_N_Mux_64_2_2_1_5072_out1 & bnn_And_64Sx64S_64S_1_5188_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5190
         assign bnn_And_64Sx64S_64S_1_5190_out1 = bnn_N_Mux_64_2_2_1_5068_out1 & bnn_And_64Sx64S_64S_1_5189_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5191
         assign bnn_And_64Sx64S_64S_1_5191_out1 = bnn_N_Mux_64_2_2_1_5064_out1 & bnn_And_64Sx64S_64S_1_5190_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5192
         assign bnn_And_64Sx64S_64S_1_5192_out1 = bnn_N_Mux_64_2_2_1_5060_out1 & bnn_And_64Sx64S_64S_1_5191_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5193
         assign bnn_And_64Sx64S_64S_1_5193_out1 = bnn_N_Mux_64_2_2_1_5056_out1 & bnn_And_64Sx64S_64S_1_5192_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5194
         assign bnn_And_64Sx64S_64S_1_5194_out1 = bnn_N_Mux_64_2_2_1_5052_out1 & bnn_And_64Sx64S_64S_1_5193_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5195
         assign bnn_And_64Sx64S_64S_1_5195_out1 = bnn_N_Mux_64_2_2_4_5048_out1 & bnn_And_64Sx64S_64S_1_5194_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5196
         assign bnn_And_64Sx64S_64S_1_5196_out1 = bnn_N_Mux_64_2_2_4_5044_out1 & bnn_And_64Sx64S_64S_1_5195_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5197
         assign bnn_And_64Sx64S_64S_1_5197_out1 = bnn_N_Mux_64_2_2_4_5040_out1 & bnn_And_64Sx64S_64S_1_5196_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5198
         assign bnn_And_64Sx64S_64S_1_5198_out1 = bnn_N_Mux_64_2_2_1_5036_out1 & bnn_And_64Sx64S_64S_1_5197_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5199
         assign bnn_And_64Sx64S_64S_1_5199_out1 = bnn_N_Mux_64_2_2_1_5032_out1 & bnn_And_64Sx64S_64S_1_5198_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5200
         assign bnn_And_64Sx64S_64S_1_5200_out1 = bnn_N_Mux_64_2_2_4_5028_out1 & bnn_And_64Sx64S_64S_1_5199_out1;

         // resource: bnn_And_64Sx64S_64S_1  instance: bnn_And_64Sx64S_64S_1_5201
         assign bnn_And_64Sx64S_64S_1_5201_out1 = bnn_N_Mux_64_2_2_1_5024_out1 & bnn_And_64Sx64S_64S_1_5200_out1;

         // resource: bnn_N_Mux_64_2_2_1
         always @(s_reg_907 or bnn_And_64Sx64S_64S_1_5201_out1)
          begin :bnn_N_Mux_64_2_2_1_5202
            if (s_reg_907) begin
               bnn_N_Mux_64_2_2_1_5202_out1 = 64'd18446744073709551615;
            end
            else begin
               bnn_N_Mux_64_2_2_1_5202_out1 = bnn_And_64Sx64S_64S_1_5201_out1;
            end
         end

         // resource: bnn_LessThan_5Ux32U_1U_4  instance: bnn_LessThan_5Ux32U_1U_4_5203
         assign bnn_LessThan_5Ux32U_1U_4_5203_out1 = {27'b000000000000000000000000000, s_reg_871} < s_reg_1000;

         // resource: bnn_LessThan_5Ux32U_1U_4  instance: bnn_LessThan_5Ux32U_1U_4_5204
         assign bnn_LessThan_5Ux32U_1U_4_5204_out1 = {27'b000000000000000000000000000, s_reg_871} < s_reg_1000;

         // resource: mux_6bx2i
         always @(bnn_Add_7Sx5S_7S_4_195_out1 or gs_ctrl599)
          begin :drive_bnn_N_Mux_12_64_13_4_5206_ctrl1
            if (gs_ctrl599) begin
               if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                  bnn_N_Mux_12_64_13_4_5206_ctrl1 = 6'd00;
               end
               else begin
                  bnn_N_Mux_12_64_13_4_5206_ctrl1 = bnn_Add_7Sx5S_7S_4_195_out1[5:0];
               end
            end
            else begin
               bnn_N_Mux_12_64_13_4_5206_ctrl1 = 6'd00;
            end
         end

         // resource: bnn_N_Mux_12_64_13_4
         always @(fixed_buffer_0_if_1_dout_wire or fixed_buffer_1_if_1_dout_wire or fixed_buffer_2_if_1_dout_wire or fixed_buffer_3_if_1_dout_wire or fixed_buffer_4_if_1_dout_wire or fixed_buffer_5_if_1_dout_wire or fixed_buffer_6_if_1_dout_wire or fixed_buffer_7_if_1_dout_wire or fixed_buffer_8_if_1_dout_wire or fixed_buffer_9_if_1_dout_wire or fixed_buffer_10_if_1_dout_wire or fixed_buffer_11_if_1_dout_wire or fixed_buffer_12_if_1_dout_wire or fixed_buffer_13_if_1_dout_wire or 
fixed_buffer_14_if_1_dout_wire
          or fixed_buffer_15_if_1_dout_wire or fixed_buffer_16_if_1_dout_wire or fixed_buffer_17_if_1_dout_wire or fixed_buffer_18_if_1_dout_wire or fixed_buffer_19_if_1_dout_wire or fixed_buffer_20_if_1_dout_wire or fixed_buffer_21_if_1_dout_wire or fixed_buffer_22_if_1_dout_wire or fixed_buffer_23_if_1_dout_wire or fixed_buffer_24_if_1_dout_wire or fixed_buffer_25_if_1_dout_wire or fixed_buffer_26_if_1_dout_wire or fixed_buffer_27_if_1_dout_wire or fixed_buffer_28_if_1_dout_wire or 
fixed_buffer_29_if_1_dout_wire
          or fixed_buffer_30_if_1_dout_wire or fixed_buffer_31_if_1_dout_wire or fixed_buffer_32_if_1_dout_wire or fixed_buffer_33_if_1_dout_wire or fixed_buffer_34_if_1_dout_wire or fixed_buffer_35_if_1_dout_wire or fixed_buffer_36_if_1_dout_wire or fixed_buffer_37_if_1_dout_wire or fixed_buffer_38_if_1_dout_wire or fixed_buffer_39_if_1_dout_wire or fixed_buffer_40_if_1_dout_wire or fixed_buffer_41_if_1_dout_wire or fixed_buffer_42_if_1_dout_wire or fixed_buffer_43_if_1_dout_wire or 
fixed_buffer_44_if_1_dout_wire
          or fixed_buffer_45_if_1_dout_wire or fixed_buffer_46_if_1_dout_wire or fixed_buffer_47_if_1_dout_wire or fixed_buffer_48_if_1_dout_wire or fixed_buffer_49_if_1_dout_wire or fixed_buffer_50_if_1_dout_wire or fixed_buffer_51_if_1_dout_wire or fixed_buffer_52_if_1_dout_wire or fixed_buffer_53_if_1_dout_wire or fixed_buffer_54_if_1_dout_wire or fixed_buffer_55_if_1_dout_wire or fixed_buffer_56_if_1_dout_wire or fixed_buffer_57_if_1_dout_wire or fixed_buffer_58_if_1_dout_wire or 
fixed_buffer_59_if_1_dout_wire
          or fixed_buffer_60_if_1_dout_wire or fixed_buffer_61_if_1_dout_wire or fixed_buffer_62_if_1_dout_wire or fixed_buffer_63_if_1_dout_wire or bnn_N_Mux_12_64_13_4_5206_ctrl1)
          begin :bnn_N_Mux_12_64_13_4_5206
            case (bnn_N_Mux_12_64_13_4_5206_ctrl1) 

               6'd01: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_1_if_1_dout_wire;
               end
               
               6'd02: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_2_if_1_dout_wire;
               end
               
               6'd03: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_3_if_1_dout_wire;
               end
               
               6'd04: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_4_if_1_dout_wire;
               end
               
               6'd05: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_5_if_1_dout_wire;
               end
               
               6'd06: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_6_if_1_dout_wire;
               end
               
               6'd07: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_7_if_1_dout_wire;
               end
               
               6'd08: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_8_if_1_dout_wire;
               end
               
               6'd09: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_9_if_1_dout_wire;
               end
               
               6'd10: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_10_if_1_dout_wire;
               end
               
               6'd11: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_11_if_1_dout_wire;
               end
               
               6'd12: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_12_if_1_dout_wire;
               end
               
               6'd13: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_13_if_1_dout_wire;
               end
               
               6'd14: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_14_if_1_dout_wire;
               end
               
               6'd15: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_15_if_1_dout_wire;
               end
               
               6'd16: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_16_if_1_dout_wire;
               end
               
               6'd17: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_17_if_1_dout_wire;
               end
               
               6'd18: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_18_if_1_dout_wire;
               end
               
               6'd19: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_19_if_1_dout_wire;
               end
               
               6'd20: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_20_if_1_dout_wire;
               end
               
               6'd21: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_21_if_1_dout_wire;
               end
               
               6'd22: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_22_if_1_dout_wire;
               end
               
               6'd23: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_23_if_1_dout_wire;
               end
               
               6'd24: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_24_if_1_dout_wire;
               end
               
               6'd25: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_25_if_1_dout_wire;
               end
               
               6'd26: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_26_if_1_dout_wire;
               end
               
               6'd27: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_27_if_1_dout_wire;
               end
               
               6'd28: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_28_if_1_dout_wire;
               end
               
               6'd29: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_29_if_1_dout_wire;
               end
               
               6'd30: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_30_if_1_dout_wire;
               end
               
               6'd31: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_31_if_1_dout_wire;
               end
               
               6'd32: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_32_if_1_dout_wire;
               end
               
               6'd33: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_33_if_1_dout_wire;
               end
               
               6'd34: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_34_if_1_dout_wire;
               end
               
               6'd35: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_35_if_1_dout_wire;
               end
               
               6'd36: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_36_if_1_dout_wire;
               end
               
               6'd37: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_37_if_1_dout_wire;
               end
               
               6'd38: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_38_if_1_dout_wire;
               end
               
               6'd39: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_39_if_1_dout_wire;
               end
               
               6'd40: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_40_if_1_dout_wire;
               end
               
               6'd41: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_41_if_1_dout_wire;
               end
               
               6'd42: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_42_if_1_dout_wire;
               end
               
               6'd43: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_43_if_1_dout_wire;
               end
               
               6'd44: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_44_if_1_dout_wire;
               end
               
               6'd45: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_45_if_1_dout_wire;
               end
               
               6'd46: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_46_if_1_dout_wire;
               end
               
               6'd47: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_47_if_1_dout_wire;
               end
               
               6'd48: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_48_if_1_dout_wire;
               end
               
               6'd49: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_49_if_1_dout_wire;
               end
               
               6'd50: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_50_if_1_dout_wire;
               end
               
               6'd51: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_51_if_1_dout_wire;
               end
               
               6'd52: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_52_if_1_dout_wire;
               end
               
               6'd53: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_53_if_1_dout_wire;
               end
               
               6'd54: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_54_if_1_dout_wire;
               end
               
               6'd55: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_55_if_1_dout_wire;
               end
               
               6'd56: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_56_if_1_dout_wire;
               end
               
               6'd57: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_57_if_1_dout_wire;
               end
               
               6'd58: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_58_if_1_dout_wire;
               end
               
               6'd59: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_59_if_1_dout_wire;
               end
               
               6'd60: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_60_if_1_dout_wire;
               end
               
               6'd61: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_61_if_1_dout_wire;
               end
               
               6'd62: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_62_if_1_dout_wire;
               end
               
               6'd63: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_63_if_1_dout_wire;
               end
               
               default: begin
                  bnn_N_Mux_12_64_13_4_5206_out1 = fixed_buffer_0_if_1_dout_wire;
               end
               
            endcase

         end

         // resource: bnn_Equal_1Ux1U_1U_1  instance: bnn_Equal_1Ux1U_1U_1_1
         assign bnn_Equal_1Ux1U_1U_1_1_out1 = !bnn_And_1Sx1U_1U_4_67_out1;

         // resource: bnn_Equal_1Ux1U_1U_1  instance: bnn_Equal_1Ux1U_1U_1_1_1
         assign bnn_Equal_1Ux1U_1U_1_1_1_out1 = !bnn_And_1Sx1U_1U_4_67_out1;

         // resource: bnn_Equal_1Ux1U_1U_1  instance: bnn_Equal_1Ux1U_1U_1_1_2
         assign bnn_Equal_1Ux1U_1U_1_1_2_out1 = !bnn_LessThan_10Ux32U_1U_4_1576_out1;

         // resource: bnn_Equal_1Ux1U_1U_1  instance: bnn_Equal_1Ux1U_1U_1_1_3
         assign bnn_Equal_1Ux1U_1U_1_1_3_out1 = !bnn_LessThan_5Ux32U_1U_4_5203_out1;

         // resource: bnn_Equal_1Ux1U_1U_1  instance: bnn_Equal_1Ux1U_1U_1_1_4
         assign bnn_Equal_1Ux1U_1U_1_1_4_out1 = !bnn_LessThan_5Ux32U_1U_4_5204_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_870_stage10
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                        end
                        else begin
                           s_reg_870_stage10 <= bnn_And_1Sx1U_1U_4_67_out1;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: regr_8b
         always @(posedge clk)
          begin :drive_s_reg_1020_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1020_stage1_slice <= bnn_Sub_8Sx2S_8S_4_1518_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1021_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1021_stage1_slice <= s_reg_1021[4:0];
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1027_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1027_stage1 <= s_reg_1027;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1029_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1029_stage1_slice <= s_reg_1029[4:0];
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1030_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1030_stage1 <= s_reg_1030;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1031_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1031_stage1_slice <= s_reg_1031[4:0];
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1032_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1032_stage1_slice <= s_reg_1032[4:0];
            end
         end

         // resource: regr_10b
         always @(posedge clk)
          begin :drive_s_reg_1034_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1034_stage1 <= s_reg_1034;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1035_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1035_stage1 <= s_reg_1035;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1036_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1036_stage1 <= s_reg_1036;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1037_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1037_stage1 <= bnn_Or_1Sx1U_1S_4_1504_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1038_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1038_stage1 <= bnn_Or_1Sx1U_1S_4_1505_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1039_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1039_stage1 <= s_reg_1039;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1040_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1040_stage1 <= bnn_GreaterThan_6Sx4S_1U_4_1506_out1;
            end
         end

         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1041_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1041_stage1_slice <= s_reg_1041[5:0];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1042_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1042_stage1 <= bnn_Or_1Sx1U_1S_4_1507_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1043_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1043_stage1 <= s_reg_1043;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1044_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1044_stage1 <= s_reg_1044;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1045_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1045_stage1 <= bnn_GreaterThan_6Sx4S_1U_4_1508_out1;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1046_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1046_stage1_slice <= s_reg_1046[4:0];
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1047_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1047_stage1 <= s_reg_1047;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1048_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1048_stage1 <= s_reg_1048;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1049_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1049_stage1 <= bnn_Or_1Sx1U_1S_4_1509_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1050_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1050_stage1 <= s_reg_1050;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1051_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1051_stage1 <= bnn_Or_1Sx1U_1S_4_1510_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1052_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1052_stage1 <= s_reg_1052;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1053_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1053_stage1 <= s_reg_1053;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1054_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1054_stage1 <= s_reg_1054;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1055_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1055_stage1 <= bnn_Or_1Sx1U_1S_4_1511_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1056_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1056_stage1 <= s_reg_1056;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1057_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1057_stage1 <= s_reg_1057;
            end
         end

         // resource: regr_6b
         always @(posedge clk)
          begin :drive_s_reg_1058_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1058_stage1_slice <= s_reg_1058[5:0];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1059_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1059_stage1 <= s_reg_1059;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1060_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1060_stage1 <= s_reg_1060;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1061_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1061_stage1 <= s_reg_1061;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1062_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1062_stage1 <= bnn_Or_1Sx1U_1S_4_1512_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1063_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1063_stage1 <= s_reg_1063;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1064_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1064_stage1 <= bnn_GreaterThan_6Sx4S_1U_4_1513_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1065_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1065_stage1 <= bnn_Or_1Sx1U_1S_4_1514_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1066_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1066_stage1 <= s_reg_1066;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1067_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1067_stage1_slice <= s_reg_1067[4:0];
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1068_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1068_stage1_slice <= s_reg_1068[4:0];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1069_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1069_stage1 <= s_reg_1068[5];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1073_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1073_stage1 <= s_reg_1073;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1074_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1074_stage1 <= s_reg_1074;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1075_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1075_stage1 <= s_reg_1075;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1076_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1076_stage1_slice <= s_reg_1076[4:0];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1079_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1079_stage1 <= s_reg_1079;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1080_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1080_stage1 <= s_reg_1080;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1081_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1081_stage1 <= s_reg_1081;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1083_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1083_stage1 <= s_reg_1083;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1085_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1085_stage1 <= s_reg_1085;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1088_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1088_stage1 <= s_reg_1088;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_1093_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1093_stage1_slice <= s_reg_1093[4:0];
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1111_stage1
            if (stall0) begin
            end
            else begin
               s_reg_1111_stage1 <= s_reg_1111;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_870_stage1
            if (stall0) begin
            end
            else begin
               s_reg_870_stage1 <= s_reg_870;
            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_s_reg_871_stage1
            if (stall0) begin
            end
            else begin
               s_reg_871_stage1 <= s_reg_871;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1044_stage10
            if (stall0) begin
            end
            else begin
               s_reg_1044_stage10 <= bnn_LessThan_5Ux32U_1U_4_5203_out1;
            end
         end

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_s_reg_1044_stage2
            if (stall0) begin
            end
            else begin
               s_reg_1044_stage2 <= s_reg_1044_stage10;
            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle1_state
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        cycle1_state <= 1'b1;
                     end
                  end
                  
                  5'd11: begin
                     if (cycle1_state) begin
                        cycle1_state <= drain2;
                     end
                     else begin
                        cycle1_state <= bnn_Equal_1Ux1U_1U_1_1_2_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle2_state
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd09: begin
                     if (!bnn_LessThan_2Ux2U_1U_4_238_out1 && (!bnn_LessThan_2Ux2U_1U_4_239_out1 && 32'd0000000000 != s_reg_1000)) begin
                        cycle2_state <= 1'b1;
                     end
                  end
                  
                  5'd11: begin
                     cycle2_state <= cycle1_state;
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         always @(vld_0 or rdy_0 or global_state)
          begin :drive_en_0
            case (global_state) 

               5'd19: begin
                  en_0 = !vld_0 | rdy_0;
               end
               
               default: begin
                  en_0 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_vld_0
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     vld_0 <= 1'b0;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        vld_0 <= 1'b0;
                     end
                  end
                  
                  5'd19: begin
                     vld_0 <= 1'b1;
                  end
                  
               endcase

            end
         end

         assign rdy_0 = (!vld_1 | rdy_1) & !iostall_1;

         // resource: mux_1bx2i
         always @(vld_0 or vld_1 or rdy_1 or iostall_1 or global_state)
          begin :drive_en_1
            case (global_state) 

               5'd19: begin
                  en_1 = (!vld_1 | rdy_1) & (!iostall_1 & vld_0);
               end
               
               default: begin
                  en_1 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_vld_1
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     vld_1 <= 1'b0;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        vld_1 <= 1'b0;
                     end
                  end
                  
                  5'd19: begin
                     vld_1 <= !iostall_1 & vld_0 | vld_1 & !rdy_1;
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         always @(iostall_2 or global_state)
          begin :drive_rdy_1
            case (global_state) 

               5'd19: begin
                  rdy_1 = !iostall_2;
               end
               
               default: begin
                  rdy_1 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(bnn_Not_1U_1U_4_10_out1 or cycle1_state2 or global_state)
          begin :drive_iostall_1
            case (global_state) 

               5'd19: begin
                  if (cycle1_state2) begin
                     iostall_1 = 1'b0;
                  end
                  else begin
                     iostall_1 = bnn_Not_1U_1U_4_10_out1;
                  end
               end
               
               default: begin
                  iostall_1 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(vld_1 or iostall_2 or global_state)
          begin :drive_en_2
            case (global_state) 

               5'd19: begin
                  en_2 = !iostall_2 & vld_1;
               end
               
               default: begin
                  en_2 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         always @(bnn_And_1Sx1U_1U_4_18_out1 or cycle2_state2 or global_state)
          begin :drive_iostall_2
            case (global_state) 

               5'd19: begin
                  case (cycle2_state2) 

                     2'd0, 2'd1: begin
                        iostall_2 = bnn_And_1Sx1U_1U_4_18_out1;
                     end
                     
                     default: begin
                        iostall_2 = 1'b0;
                     end
                     
                  endcase

               end
               
               default: begin
                  iostall_2 = 1'b0;
               end
               
            endcase

         end

         // resource: mux_1bx4i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle1_state2
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     cycle1_state2 <= 1'b1;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        cycle1_state2 <= 1'b1;
                     end
                  end
                  
                  5'd19: begin
                     if (en_0) begin
                        if (en_1) begin
                           if (cycle1_state2) begin
                              cycle1_state2 <= drain3;
                           end
                           else begin
                              case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                                 7'd001: begin
                                    cycle1_state2 <= bnn_Equal_1Ux1U_1U_1_1_1_out1;
                                 end
                                 
                                 default: begin
                                    cycle1_state2 <= bnn_Equal_1Ux1U_1U_1_1_out1;
                                 end
                                 
                              endcase

                           end
                        end
                        else begin
                           cycle1_state2 <= drain3;
                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_cycle2_state2
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd00: begin
                     cycle2_state2 <= 2'd2;
                  end
                  
                  5'd18: begin
                     if (bnn_Add_7Sx5S_7S_4_195_out1[6] && s_reg_907) begin
                        cycle2_state2 <= 2'd2;
                     end
                  end
                  
                  5'd19: begin
                     if (en_1) begin
                        if (cycle1_state2) begin
                           cycle2_state2 <= 2'd2;
                        end
                        else begin
                           case (bnn_N_MuxB_160_2_0_4_37_out1[159:153]) 

                              7'd001: begin
                                 cycle2_state2 <= 2'd0;
                              end
                              
                              default: begin
                                 cycle2_state2 <= 2'd1;
                              end
                              
                           endcase

                        end
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle1_state0
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        cycle1_state0 <= 1'b1;
                     end
                  end
                  
                  5'd15: begin
                     if (cycle1_state0) begin
                        cycle1_state0 <= drain1;
                     end
                     else begin
                        cycle1_state0 <= bnn_Equal_1Ux1U_1U_1_1_3_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle2_state0
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        cycle2_state0 <= 1'b1;
                     end
                  end
                  
                  5'd15: begin
                     cycle2_state0 <= cycle1_state0;
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle3_state
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        cycle3_state <= 1'b1;
                     end
                  end
                  
                  5'd15: begin
                     cycle3_state <= cycle2_state0;
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx3i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle1_state1
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (!s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        cycle1_state1 <= 1'b1;
                     end
                  end
                  
                  5'd16: begin
                     if (cycle1_state1) begin
                        cycle1_state1 <= drain;
                     end
                     else begin
                        cycle1_state1 <= bnn_Equal_1Ux1U_1U_1_1_4_out1;
                     end
                  end
                  
               endcase

            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_cycle2_state1
            if (stall0) begin
            end
            else begin
               case (global_state) 

                  5'd14: begin
                     if (!s_reg_1006 && 32'd0000000000 != s_reg_1000) begin
                        cycle2_state1 <= 1'b1;
                     end
                  end
                  
                  5'd16: begin
                     cycle2_state1 <= cycle1_state1;
                  end
                  
               endcase

            end
         end

         // resource: regr_5b
         always @(posedge clk)
          begin :drive_global_state
            if (reset == 1'b1) begin
               global_state <= 5'd00;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  global_state <= global_state_next;
               end
            end
         end

         // resource: mux_5bx14i
         always @(s_reg_1000 or s_reg_1005[31:0] or s_reg_1006 or s_reg_1112 or s_reg_907 or bnn_Add_5Sx4S_6S_1_180_out1[4] or bnn_Add_7Sx5S_7S_4_195_out1[6] or bnn_LessThan_2Ux2U_1U_4_238_out1 or bnn_LessThan_2Ux2U_1U_4_239_out1 or bnn_LessThan_10Ux32U_1U_4_4104_out1 or bnn_N_Mux_3_2_6_4_4105_out1 or s_reg_870_stage10 or s_reg_1044_stage2 or cycle2_state or en_2 or cycle2_state2 or cycle3_state or cycle2_state1 or global_state)
          begin :drive_global_state_next
            case (global_state) 

               5'd00: begin
                  global_state_next = 5'd19;
               end
               
               5'd01, 5'd02: begin
                  if (bnn_Add_5Sx4S_6S_1_180_out1[4]) begin
                     case (s_reg_1005[31:0]) 

                        32'd0000000000: begin
                           global_state_next = 5'd03;
                        end
                        
                        default: begin
                           global_state_next = 5'd07;
                        end
                        
                     endcase

                  end
                  else begin
                     global_state_next = 5'd02;
                  end
               end
               
               5'd04: begin
                  global_state_next = 5'd13;
               end
               
               5'd06, 5'd08, 5'd10: begin
                  global_state_next = 5'd09;
               end
               
               5'd09: begin
                  if (bnn_LessThan_2Ux2U_1U_4_238_out1) begin
                     global_state_next = global_state + 5'd01;
                  end
                  else begin
                     if (bnn_LessThan_2Ux2U_1U_4_239_out1) begin
                        global_state_next = 5'd09;
                     end
                     else begin
                        /* state45 */
                        case (s_reg_1000) 

                           32'd0000000000: begin
                              global_state_next = 5'd12;
                           end
                           
                           default: begin
                              global_state_next = 5'd11;
                           end
                           
                        endcase

                     end
                  end
               end
               
               5'd11: begin
                  if (!cycle2_state && !s_reg_1112) begin
                     global_state_next = global_state + 5'd01;
                  end
                  else begin
                     global_state_next = 5'd11;
                  end
               end
               
               5'd12: begin
                  if (bnn_LessThan_10Ux32U_1U_4_4104_out1) begin
                     case (bnn_N_Mux_3_2_6_4_4105_out1) 

                        3'd0: begin
                           global_state_next = 5'd07;
                        end
                        
                        default: begin
                           global_state_next = 5'd05;
                        end
                        
                     endcase

                  end
                  else begin
                     global_state_next = global_state + 5'd01;
                  end
               end
               
               5'd14: begin
                  if (s_reg_1006) begin
                     case (s_reg_1000) 

                        32'd0000000000: begin
                           global_state_next = 5'd17;
                        end
                        
                        default: begin
                           global_state_next = global_state + 5'd01;
                        end
                        
                     endcase

                  end
                  else begin
                     case (s_reg_1000) 

                        32'd0000000000: begin
                           global_state_next = 5'd17;
                        end
                        
                        default: begin
                           global_state_next = 5'd16;
                        end
                        
                     endcase

                  end
               end
               
               5'd15: begin
                  if (!cycle3_state && !s_reg_1044_stage2) begin
                     global_state_next = 5'd17;
                  end
                  else begin
                     global_state_next = 5'd15;
                  end
               end
               
               5'd16: begin
                  if (!cycle2_state1 && !s_reg_907) begin
                     global_state_next = global_state + 5'd01;
                  end
                  else begin
                     global_state_next = 5'd16;
                  end
               end
               
               5'd18: begin
                  if (bnn_Add_7Sx5S_7S_4_195_out1[6]) begin
                     if (s_reg_907) begin
                        global_state_next = global_state + 5'd01;
                     end
                     else begin
                        global_state_next = 5'd17;
                     end
                  end
                  else begin
                     global_state_next = 5'd17;
                  end
               end
               
               5'd19: begin
                  if (en_2) begin
                     case (cycle2_state2) 

                        2'd0, 2'd1: begin
                           if (s_reg_870_stage10) begin
                              global_state_next = 5'd19;
                           end
                           else begin
                              global_state_next = 5'd01;
                           end
                        end
                        
                        default: begin
                           global_state_next = 5'd19;
                        end
                        
                     endcase

                  end
                  else begin
                     global_state_next = 5'd19;
                  end
               end
               
               default: begin
                  global_state_next = global_state + 5'd01;
               end
               
            endcase

         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl0
            if (reset == 1'b1) begin
               gs_ctrl0 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd15, 5'd16: begin
                        gs_ctrl0 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl0 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl4
            if (reset == 1'b1) begin
               gs_ctrl4 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd19: begin
                        gs_ctrl4 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl4 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl23
            if (reset == 1'b1) begin
               gs_ctrl23 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd12: begin
                        gs_ctrl23 <= 2'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl23 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl23 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl61
            if (reset == 1'b1) begin
               gs_ctrl61 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd15: begin
                        gs_ctrl61 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl61 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl74
            if (reset == 1'b1) begin
               gs_ctrl74 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd12: begin
                        gs_ctrl74 <= 2'd1;
                     end
                     
                     5'd15, 5'd16: begin
                        gs_ctrl74 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl74 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl105
            if (reset == 1'b1) begin
               gs_ctrl105 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd12: begin
                        gs_ctrl105 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl105 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl196
            if (reset == 1'b1) begin
               gs_ctrl196 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11: begin
                        gs_ctrl196 <= 2'd1;
                     end
                     
                     5'd12: begin
                        gs_ctrl196 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl196 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl197
            if (reset == 1'b1) begin
               gs_ctrl197 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11: begin
                        gs_ctrl197 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl197 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl198
            if (reset == 1'b1) begin
               gs_ctrl198 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11, 5'd19: begin
                        gs_ctrl198 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl198 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl199
            if (reset == 1'b1) begin
               gs_ctrl199 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11: begin
                        gs_ctrl199 <= 2'd1;
                     end
                     
                     5'd19: begin
                        gs_ctrl199 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl199 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx6i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl205
            if (reset == 1'b1) begin
               gs_ctrl205 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd02, 5'd17: begin
                        gs_ctrl205 <= 3'd1;
                     end
                     
                     5'd06, 5'd08: begin
                        gs_ctrl205 <= 3'd2;
                     end
                     
                     5'd09: begin
                        gs_ctrl205 <= 3'd3;
                     end
                     
                     5'd10: begin
                        gs_ctrl205 <= 3'd4;
                     end
                     
                     5'd11: begin
                        gs_ctrl205 <= 3'd5;
                     end
                     
                     default: begin
                        gs_ctrl205 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx5i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl206
            if (reset == 1'b1) begin
               gs_ctrl206 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd06, 5'd08: begin
                        gs_ctrl206 <= 3'd1;
                     end
                     
                     5'd09: begin
                        gs_ctrl206 <= 3'd2;
                     end
                     
                     5'd10: begin
                        gs_ctrl206 <= 3'd3;
                     end
                     
                     5'd11: begin
                        gs_ctrl206 <= 3'd4;
                     end
                     
                     default: begin
                        gs_ctrl206 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx5i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl210
            if (reset == 1'b1) begin
               gs_ctrl210 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd06, 5'd08: begin
                        gs_ctrl210 <= 3'd1;
                     end
                     
                     5'd09: begin
                        gs_ctrl210 <= 3'd2;
                     end
                     
                     5'd11: begin
                        gs_ctrl210 <= 3'd3;
                     end
                     
                     5'd15, 5'd16: begin
                        gs_ctrl210 <= 3'd4;
                     end
                     
                     default: begin
                        gs_ctrl210 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl211
            if (reset == 1'b1) begin
               gs_ctrl211 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd06, 5'd08, 5'd09: begin
                        gs_ctrl211 <= 2'd1;
                     end
                     
                     5'd11: begin
                        gs_ctrl211 <= 2'd2;
                     end
                     
                     5'd15, 5'd16: begin
                        gs_ctrl211 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl211 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx6i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl214
            if (reset == 1'b1) begin
               gs_ctrl214 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd06, 5'd08: begin
                        gs_ctrl214 <= 3'd1;
                     end
                     
                     5'd09: begin
                        gs_ctrl214 <= 3'd2;
                     end
                     
                     5'd10: begin
                        gs_ctrl214 <= 3'd3;
                     end
                     
                     5'd11: begin
                        gs_ctrl214 <= 3'd4;
                     end
                     
                     5'd15, 5'd16: begin
                        gs_ctrl214 <= 3'd5;
                     end
                     
                     default: begin
                        gs_ctrl214 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl217
            if (reset == 1'b1) begin
               gs_ctrl217 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd09: begin
                        gs_ctrl217 <= 2'd1;
                     end
                     
                     5'd11: begin
                        gs_ctrl217 <= 2'd2;
                     end
                     
                     5'd18: begin
                        gs_ctrl217 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl217 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl219
            if (reset == 1'b1) begin
               gs_ctrl219 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11, 5'd12: begin
                        gs_ctrl219 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl219 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl222
            if (reset == 1'b1) begin
               gs_ctrl222 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd10: begin
                        gs_ctrl222 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl222 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl224
            if (reset == 1'b1) begin
               gs_ctrl224 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd10: begin
                        gs_ctrl224 <= 2'd1;
                     end
                     
                     5'd11: begin
                        gs_ctrl224 <= 2'd2;
                     end
                     
                     5'd12: begin
                        gs_ctrl224 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl224 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl226
            if (reset == 1'b1) begin
               gs_ctrl226 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd10: begin
                        gs_ctrl226 <= 2'd1;
                     end
                     
                     5'd11: begin
                        gs_ctrl226 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl226 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl228
            if (reset == 1'b1) begin
               gs_ctrl228 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd09: begin
                        gs_ctrl228 <= 2'd1;
                     end
                     
                     5'd10: begin
                        gs_ctrl228 <= 2'd2;
                     end
                     
                     5'd11: begin
                        gs_ctrl228 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl228 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl240
            if (reset == 1'b1) begin
               gs_ctrl240 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd08: begin
                        gs_ctrl240 <= 2'd1;
                     end
                     
                     5'd11: begin
                        gs_ctrl240 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl240 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl242
            if (reset == 1'b1) begin
               gs_ctrl242 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd11: begin
                        gs_ctrl242 <= 2'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl242 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl242 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl264
            if (reset == 1'b1) begin
               gs_ctrl264 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd12: begin
                        gs_ctrl264 <= 2'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl264 <= 2'd2;
                     end
                     
                     5'd16: begin
                        gs_ctrl264 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl264 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx3i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl266
            if (reset == 1'b1) begin
               gs_ctrl266 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd14, 5'd16, 5'd18: begin
                        gs_ctrl266 <= 2'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl266 <= 2'd2;
                     end
                     
                     default: begin
                        gs_ctrl266 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_2bx4i
         // resource: regr_2b
         always @(posedge clk)
          begin :drive_gs_ctrl267
            if (reset == 1'b1) begin
               gs_ctrl267 <= 2'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd14, 5'd16: begin
                        gs_ctrl267 <= 2'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl267 <= 2'd2;
                     end
                     
                     5'd18: begin
                        gs_ctrl267 <= 2'd3;
                     end
                     
                     default: begin
                        gs_ctrl267 <= 2'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl599
            if (reset == 1'b1) begin
               gs_ctrl599 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd18: begin
                        gs_ctrl599 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl599 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl690
            if (reset == 1'b1) begin
               gs_ctrl690 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd01, 5'd02: begin
                        gs_ctrl690 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl690 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_1bx2i
         // resource: regr_1b
         always @(posedge clk)
          begin :drive_gs_ctrl691
            if (reset == 1'b1) begin
               gs_ctrl691 <= 1'b0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd02: begin
                        gs_ctrl691 <= 1'b1;
                     end
                     
                     default: begin
                        gs_ctrl691 <= 1'b0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx5i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl692
            if (reset == 1'b1) begin
               gs_ctrl692 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd14: begin
                        gs_ctrl692 <= 3'd1;
                     end
                     
                     5'd15: begin
                        gs_ctrl692 <= 3'd2;
                     end
                     
                     5'd16: begin
                        gs_ctrl692 <= 3'd3;
                     end
                     
                     5'd18: begin
                        gs_ctrl692 <= 3'd4;
                     end
                     
                     default: begin
                        gs_ctrl692 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         // resource: mux_3bx6i
         // resource: regr_3b
         always @(posedge clk)
          begin :drive_gs_ctrl820
            if (reset == 1'b1) begin
               gs_ctrl820 <= 3'd0;
            end
            else begin
               if (stall0) begin
               end
               else begin
                  case (global_state_next) 

                     5'd12: begin
                        gs_ctrl820 <= 3'd1;
                     end
                     
                     5'd14: begin
                        gs_ctrl820 <= 3'd2;
                     end
                     
                     5'd15: begin
                        gs_ctrl820 <= 3'd3;
                     end
                     
                     5'd16: begin
                        gs_ctrl820 <= 3'd4;
                     end
                     
                     5'd18: begin
                        gs_ctrl820 <= 3'd5;
                     end
                     
                     default: begin
                        gs_ctrl820 <= 3'd0;
                     end
                     
                  endcase

               end
            end
         end

         assign xcelreq_busy = bnn_Or_1Sx1U_1S_4_6_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_3
         assign bnn_Or_1Sx1U_1S_4_3_out1 = xcelreq_m_unvalidated_req | xcelreq_vld;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_4
         assign bnn_And_1Sx1U_1U_4_4_out1 = bnn_Or_1Sx1U_1S_4_3_out1 & xcelreq_m_busy_req_0;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_6
         assign bnn_Or_1Sx1U_1S_4_6_out1 = bnn_And_1Sx1U_1U_4_4_out1 | xcelreq_m_stall_reg_full;

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_7
         assign bnn_Not_1U_1U_4_7_out1 = !bnn_Or_1Sx1U_1S_4_6_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_8
         assign bnn_And_1Sx1U_1U_4_8_out1 = bnn_Not_1U_1U_4_7_out1 & xcelreq_vld;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_9
         assign bnn_Or_1Sx1U_1S_4_9_out1 = bnn_And_1Sx1U_1U_4_8_out1 | xcelreq_m_stall_reg_full;

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_10
         assign bnn_Not_1U_1U_4_10_out1 = !bnn_Or_1Sx1U_1S_4_9_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelreq_m_unvalidated_req
            if (reset == 1'b1) begin
               xcelreq_m_unvalidated_req <= 1'd1;
            end
            else begin
               xcelreq_m_unvalidated_req <= bnn_N_Muxb_1_2_18_4_1_out1;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(xcelreq_vld or xcelreq_m_busy_req_0 or xcelreq_m_unvalidated_req)
          begin :bnn_N_Muxb_1_2_18_4_1
            if (xcelreq_m_busy_req_0) begin
               bnn_N_Muxb_1_2_18_4_1_out1 = xcelreq_m_unvalidated_req;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_1_out1 = xcelreq_vld;
            end
         end

         // resource: regr_160b
         always @(posedge clk)
          begin :drive_xcelreq_m_stall_reg
            if (bnn_And_1Sx1U_1U_4_13_out1) begin
               xcelreq_m_stall_reg <= xcelreq_data;
            end
         end

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_11
         assign bnn_Not_1U_1U_4_11_out1 = !xcelreq_m_stall_reg_full;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_12
         assign bnn_And_1Sx1U_1U_4_12_out1 = bnn_Or_1Sx1U_1S_4_9_out1 & xcelreq_m_stalling;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_13
         assign bnn_And_1Sx1U_1U_4_13_out1 = bnn_And_1Sx1U_1U_4_12_out1 & bnn_Not_1U_1U_4_11_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelreq_m_stall_reg_full
            if (reset == 1'b1) begin
               xcelreq_m_stall_reg_full <= 1'd0;
            end
            else begin
               xcelreq_m_stall_reg_full <= bnn_And_1Sx1U_1U_4_14_out1;
            end
         end

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_14
         assign bnn_And_1Sx1U_1U_4_14_out1 = bnn_Or_1Sx1U_1S_4_9_out1 & xcelreq_m_stalling;

         assign xcelresp_vld = bnn_Or_1Sx1U_1S_4_17_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_17
         assign bnn_Or_1Sx1U_1S_4_17_out1 = xcelresp_m_unacked_req | bnn_Xor_1Ux1U_1U_4_16_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelresp_m_unacked_req
            if (reset == 1'b1) begin
               xcelresp_m_unacked_req <= 1'd0;
            end
            else begin
               xcelresp_m_unacked_req <= bnn_And_1Sx1U_1U_4_18_out1;
            end
         end

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_18
         assign bnn_And_1Sx1U_1U_4_18_out1 = xcelresp_busy & xcelresp_vld;

         // resource: bnn_Xor_1Ux1U_1U_4  instance: bnn_Xor_1Ux1U_1U_4_16
         assign bnn_Xor_1Ux1U_1U_4_16_out1 = xcelresp_m_req_m_trig_req ^ xcelresp_m_req_m_prev_trig_req;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_xcelresp_m_req_m_prev_trig_req
            if (reset == 1'b1) begin
               xcelresp_m_req_m_prev_trig_req <= 1'd0;
            end
            else begin
               xcelresp_m_req_m_prev_trig_req <= xcelresp_m_req_m_trig_req;
            end
         end

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_19
         assign bnn_Not_1U_1U_4_19_out1 = !xcelresp_m_req_m_trig_req;

         assign memreq_vld = bnn_Or_1Sx1U_1S_4_21_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_21
         assign bnn_Or_1Sx1U_1S_4_21_out1 = memreq_m_unacked_req | bnn_Xor_1Ux1U_1U_4_20_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memreq_m_unacked_req
            if (reset == 1'b1) begin
               memreq_m_unacked_req <= 1'd0;
            end
            else begin
               memreq_m_unacked_req <= bnn_And_1Sx1U_1U_4_22_out1;
            end
         end

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_22
         assign bnn_And_1Sx1U_1U_4_22_out1 = memreq_busy & memreq_vld;

         // resource: bnn_Xor_1Ux1U_1U_4  instance: bnn_Xor_1Ux1U_1U_4_20
         assign bnn_Xor_1Ux1U_1U_4_20_out1 = memreq_m_req_m_trig_req ^ memreq_m_req_m_prev_trig_req;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memreq_m_req_m_prev_trig_req
            if (reset == 1'b1) begin
               memreq_m_req_m_prev_trig_req <= 1'd0;
            end
            else begin
               memreq_m_req_m_prev_trig_req <= memreq_m_req_m_trig_req;
            end
         end

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_23
         assign bnn_Not_1U_1U_4_23_out1 = !memreq_m_req_m_trig_req;

         assign memresp_busy = bnn_Or_1Sx1U_1S_4_27_out1;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_24
         assign bnn_Or_1Sx1U_1S_4_24_out1 = memresp_m_unvalidated_req | memresp_vld;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_25
         assign bnn_And_1Sx1U_1U_4_25_out1 = bnn_Or_1Sx1U_1S_4_24_out1 & memresp_m_busy_req_0;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_27
         assign bnn_Or_1Sx1U_1S_4_27_out1 = bnn_And_1Sx1U_1U_4_25_out1 | memresp_m_stall_reg_full;

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_28
         assign bnn_Not_1U_1U_4_28_out1 = !bnn_Or_1Sx1U_1S_4_27_out1;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_29
         assign bnn_And_1Sx1U_1U_4_29_out1 = bnn_Not_1U_1U_4_28_out1 & memresp_vld;

         // resource: bnn_Or_1Sx1U_1S_4  instance: bnn_Or_1Sx1U_1S_4_30
         assign bnn_Or_1Sx1U_1S_4_30_out1 = bnn_And_1Sx1U_1U_4_29_out1 | memresp_m_stall_reg_full;

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_31
         assign bnn_Not_1U_1U_4_31_out1 = !bnn_Or_1Sx1U_1S_4_30_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memresp_m_unvalidated_req
            if (reset == 1'b1) begin
               memresp_m_unvalidated_req <= 1'd1;
            end
            else begin
               memresp_m_unvalidated_req <= bnn_N_Muxb_1_2_18_4_2_out1;
            end
         end

         // resource: bnn_N_Muxb_1_2_18_4
         always @(memresp_vld or memresp_m_busy_req_0 or memresp_m_unvalidated_req)
          begin :bnn_N_Muxb_1_2_18_4_2
            if (memresp_m_busy_req_0) begin
               bnn_N_Muxb_1_2_18_4_2_out1 = memresp_m_unvalidated_req;
            end
            else begin
               bnn_N_Muxb_1_2_18_4_2_out1 = memresp_vld;
            end
         end

         // resource: regr_64b
         always @(posedge clk)
          begin :drive_memresp_m_stall_reg
            if (bnn_And_1Sx1U_1U_4_34_out1) begin
               memresp_m_stall_reg_slice <= memresp_data[63:0];
            end
         end

         // resource: bnn_Not_1U_1U_4  instance: bnn_Not_1U_1U_4_32
         assign bnn_Not_1U_1U_4_32_out1 = !memresp_m_stall_reg_full;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_33
         assign bnn_And_1Sx1U_1U_4_33_out1 = bnn_Or_1Sx1U_1S_4_30_out1 & stall0;

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_34
         assign bnn_And_1Sx1U_1U_4_34_out1 = bnn_And_1Sx1U_1U_4_33_out1 & bnn_Not_1U_1U_4_32_out1;

         // resource: regr_1b
         always @(posedge clk)
          begin :drive_memresp_m_stall_reg_full
            if (reset == 1'b1) begin
               memresp_m_stall_reg_full <= 1'd0;
            end
            else begin
               memresp_m_stall_reg_full <= bnn_And_1Sx1U_1U_4_35_out1;
            end
         end

         // resource: bnn_And_1Sx1U_1U_4  instance: bnn_And_1Sx1U_1U_4_35
         assign bnn_And_1Sx1U_1U_4_35_out1 = bnn_Or_1Sx1U_1S_4_30_out1 & stall0;

         assign memreq_data = {{2'b00, memreq_data_slice[96]}, {8'd000, {memreq_data_slice[95:64], {3'd0, memreq_data_slice[63:0]}}}};


endmodule

`timescale 1ps / 1ps
module bnn_Mod_6Ux32U_7U_4(
          in2,
          in1,
          out1,
          clk,
          stall
);
   input [5:0] in2;
   input [31:0] in1;
   output [6:0] out1;
   input clk;
   input stall;
wire in2_2, sub_115_2_n_1, sub_115_2_n_10, sub_115_2_n_12, sub_115_2_n_13,
     sub_115_2_n_14, sub_115_2_n_16, sub_115_2_n_17, sub_115_2_n_19,
     sub_115_2_n_2, sub_115_2_n_20, sub_115_2_n_21, sub_115_2_n_23,
     sub_115_2_n_24, sub_115_2_n_25, sub_115_2_n_3, sub_115_2_n_4, sub_115_2_n_5,
     sub_115_2_n_6, sub_115_2_n_7, sub_115_2_n_8, sub_115_2_n_9, sub_134_2_n_0,
     sub_134_2_n_10, sub_134_2_n_11, sub_134_2_n_12, sub_134_2_n_13,
     sub_134_2_n_14, sub_134_2_n_15, sub_134_2_n_17, sub_134_2_n_18,
     sub_134_2_n_19, sub_134_2_n_2, sub_134_2_n_20, sub_134_2_n_22,
     sub_134_2_n_23, sub_134_2_n_24, sub_134_2_n_28, sub_134_2_n_29,
     sub_134_2_n_3, sub_134_2_n_31, sub_134_2_n_4, sub_134_2_n_5, sub_134_2_n_6,
     sub_134_2_n_7, sub_134_2_n_8, sub_134_2_n_9, sub_153_2_n_0, sub_153_2_n_10,
     sub_153_2_n_11, sub_153_2_n_12, sub_153_2_n_13, sub_153_2_n_14,
     sub_153_2_n_15, sub_153_2_n_16, sub_153_2_n_19, sub_153_2_n_2,
     sub_153_2_n_20, sub_153_2_n_21, sub_153_2_n_22, sub_153_2_n_23,
     sub_153_2_n_24, sub_153_2_n_26, sub_153_2_n_27, sub_153_2_n_28,
     sub_153_2_n_3, sub_153_2_n_32, sub_153_2_n_35, sub_153_2_n_5, sub_153_2_n_7,
     sub_153_2_n_8, sub_153_2_n_9, sub_58_2_n_1, sub_58_2_n_10, sub_58_2_n_11,
     sub_58_2_n_12, sub_58_2_n_3, sub_58_2_n_4, sub_58_2_n_5, sub_58_2_n_6,
     sub_58_2_n_7, sub_58_2_n_8, sub_58_2_n_9, sub_77_2_n_1, sub_77_2_n_11,
     sub_77_2_n_12, sub_77_2_n_13, sub_77_2_n_14, sub_77_2_n_15, sub_77_2_n_16,
     sub_77_2_n_17, sub_77_2_n_2, sub_77_2_n_3, sub_77_2_n_4, sub_77_2_n_5,
     sub_77_2_n_6, sub_77_2_n_7, sub_77_2_n_9, sub_96_2_n_1, sub_96_2_n_10,
     sub_96_2_n_11, sub_96_2_n_13, sub_96_2_n_14, sub_96_2_n_16, sub_96_2_n_17,
     sub_96_2_n_18, sub_96_2_n_19, sub_96_2_n_2, sub_96_2_n_20, sub_96_2_n_3,
     sub_96_2_n_4, sub_96_2_n_5, sub_96_2_n_6, sub_96_2_n_7, sub_96_2_n_8, clk,
     stall, n_7, n_9, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20,
     n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32,
     n_33, n_34, n_35, n_36, n_37, n_38, n_40, n_42, n_43, n_72, n_73, n_74,
     n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_87, n_88,
     n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_98, n_99, n_100, n_101,
     n_104, in2_10_0_, in2_10_1_, in2_10_2_, in2_10_32_, in2_10_3_, in2_11_0_,
     in2_11_1_, in2_11_2_, in2_11_3_, in2_14_0_, in2_14_1_, in2_14_2_, in2_14_3_,
     in2_14_4_, in2_16_1_, in2_16_2_, in2_16_32_, in2_16_3_, in2_16_4_,
     in2_16_5_, in2_1_0_, in2_1_32_, in2_4_0_, in2_4_1_, in2_4_32_, in2_5_0_,
     in2_5_1_, in2_7_0_, in2_7_1_, in2_7_2_, in2_7_32_, in2_8_0_, in2_8_1_,
     in2_8_2_;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_10_reg_reg_IQ <= n_42;
 assign n_82 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 wire retime_s1_11_reg_reg_IQN;
 assign retime_s1_11_reg_reg_IQN = !retime_s1_11_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_11_reg_reg_IQ <= n_43;
 assign n_83 = retime_s1_11_reg_reg_IQN;
 reg retime_s1_12_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_12_reg_reg_IQ <= n_31;
 assign n_84 = retime_s1_12_reg_reg_IQ;
 reg retime_s1_13_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_13_reg_reg_IQ <= n_35;
 assign n_85 = retime_s1_13_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_14_reg_reg_IQ <= {in1[1]};
 assign n_87 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_15_reg_reg_IQ <= n_25;
 assign n_88 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_16_reg_reg_IQ <= {in1[2]};
 assign n_89 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_17_reg_reg_IQ <= {in1[5]};
 assign n_90 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_18_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_18_reg_reg_IQ <= {in1[15]};
 assign n_91 = retime_s1_18_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_19_reg_reg_IQ <= {in2[1]};
 assign n_92 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_1_reg_reg_IQ <= in2_11_2_;
 assign n_72 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_20_reg_reg_IQ <= {in1[14]};
 assign n_93 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 wire retime_s1_21_reg_reg_IQN;
 assign retime_s1_21_reg_reg_IQN = !retime_s1_21_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_21_reg_reg_IQ <= n_15;
 assign n_94 = retime_s1_21_reg_reg_IQN;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_22_reg_reg_IQ <= in2_11_0_;
 assign n_95 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_23_reg_reg_IQ <= {in1[13]};
 assign n_96 = retime_s1_23_reg_reg_IQ;
 reg retime_s1_24_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_24_reg_reg_IQ <= {in1[12]};
 assign n_98 = retime_s1_24_reg_reg_IQ;
 reg retime_s1_25_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_25_reg_reg_IQ <= {in1[4]};
 assign n_99 = retime_s1_25_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_26_reg_reg_IQ <= {in1[3]};
 assign n_100 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_27_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_27_reg_reg_IQ <= {in2[0]};
 assign n_101 = retime_s1_27_reg_reg_IQ;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_2_reg_reg_IQ <= n_26;
 assign n_73 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_3_reg_reg_IQ <= n_27;
 assign n_74 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 wire retime_s1_4_reg_reg_IQN;
 assign retime_s1_4_reg_reg_IQN = !retime_s1_4_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_4_reg_reg_IQ <= n_14;
 assign n_76 = retime_s1_4_reg_reg_IQN;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_5_reg_reg_IQ <= n_30;
 assign n_77 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_6_reg_reg_IQ;
 wire retime_s1_6_reg_reg_IQN;
 assign retime_s1_6_reg_reg_IQN = !retime_s1_6_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_6_reg_reg_IQ <= n_16;
 assign n_78 = retime_s1_6_reg_reg_IQN;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_7_reg_reg_IQ <= in2_11_1_;
 assign n_79 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 wire retime_s1_8_reg_reg_IQN;
 assign retime_s1_8_reg_reg_IQN = !retime_s1_8_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_8_reg_reg_IQ <= n_104;
 assign n_80 = retime_s1_8_reg_reg_IQN;
 reg retime_s1_9_reg_reg_IQ;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_9_reg_reg_IQ <= in2_11_3_;
 assign n_81 = retime_s1_9_reg_reg_IQ;
 assign {out1[0]} = ((n_82 & ~in2_16_32_) | (n_101 & in2_16_32_));
 assign in2_16_32_ = ~((n_23 & n_32) & (sub_153_2_n_24 | n_7));
 assign sub_153_2_n_26 = ~(sub_153_2_n_8 | (n_83 & sub_153_2_n_7));
 assign n_7 = ~((~sub_153_2_n_3 | sub_153_2_n_14) | sub_153_2_n_32);
 assign sub_153_2_n_8 = ~(n_87 | ~in2_14_0_);
 assign sub_153_2_n_7 = ~(~in2_14_0_ & n_87);
 assign sub_153_2_n_14 = ~(~n_99 | in2_14_3_);
 assign sub_153_2_n_3 = ~(~in2_14_4_ & n_90);
 assign sub_153_2_n_10 = ~(~n_89 & in2_14_1_);
 assign sub_153_2_n_9 = ~(~n_89 | in2_14_1_);
 assign sub_153_2_n_5 = ~(~n_90 & in2_14_4_);
 assign sub_153_2_n_2 = ~(~n_99 & in2_14_3_);
 assign sub_153_2_n_13 = ~(n_100 | ~in2_14_2_);
 assign sub_153_2_n_11 = ~(~in2_14_2_ & n_100);
 assign n_42 = ~((~stall | ~n_82) & (stall | n_17));
 assign n_43 = ~((~stall & ~n_18) | (stall & n_83));
 assign n_14 = ~(n_28 | (stall & n_76));
 assign n_16 = ~(n_29 | (stall & n_78));
 assign in2_14_0_ = ((n_84 & ~n_9) | (n_92 & n_9));
 assign in2_14_4_ = ((n_74 & ~n_9) | (n_81 & n_9));
 assign in2_14_1_ = ((n_85 & ~n_9) | (n_95 & n_9));
 assign in2_14_2_ = ((n_80 & ~n_9) | (n_79 & n_9));
 assign in2_14_3_ = ~((~n_72 | ~n_9) & (n_73 | n_9));
 assign n_28 = ~((({in1[23]} | stall) | {in1[22]}) | sub_153_2_n_28);
 assign n_29 = ~((({in1[19]} | stall) | {in1[18]}) | sub_134_2_n_24);
 assign n_15 = ~(n_33 | (stall & n_94));
 assign n_30 = ~(((sub_134_2_n_15 & sub_134_2_n_31) & ~{in1[14]}) & ~{in1[15]});
 assign n_18 = (n_40 & {in1[0]});
 assign n_17 = (n_40 ^ {in1[0]});
 assign n_31 = ~(sub_134_2_n_4 & (~{in2[1]} | {in1[0]}));
 assign n_9 = ~((~n_77 & n_78) & n_24);
 assign n_33 = ~(({in1[7]} | stall) | {in1[6]});
 assign n_32 = ~((n_91 | ~n_76) | ~n_88);
 assign n_23 = ~((n_93 | ~n_94) | ~n_24);
 assign in2_11_1_ = ~(n_19 & (~in2_10_1_ | n_37));
 assign in2_11_0_ = ~(n_36 & (~in2_10_0_ | in2_10_32_));
 assign in2_11_2_ = ~(n_11 & (~in2_10_2_ | n_20));
 assign in2_11_3_ = ~(n_12 & (~in2_10_3_ | n_13));
 assign n_34 = ~(sub_134_2_n_18 ^ sub_134_2_n_22);
 assign n_35 = ~(sub_134_2_n_4 ^ sub_134_2_n_17);
 assign n_25 = ~((({in1[9]} | {in1[10]}) | {in1[11]}) | {in1[8]});
 assign in2_16_1_ = ~(sub_153_2_n_21 ^ n_83);
 assign n_26 = (sub_134_2_n_19 ^ sub_134_2_n_0);
 assign n_27 = ~(sub_134_2_n_20 ^ sub_134_2_n_28);
 assign n_11 = ~(in2_8_1_ & n_21);
 assign n_36 = ~({in2[2]} & in2_10_32_);
 assign n_19 = ~(in2_8_0_ & n_20);
 assign n_12 = ~(in2_8_2_ & n_13);
 assign n_24 = ~(n_98 | n_96);
 assign n_40 = ~{in2[0]};
 assign n_37 = ~n_38;
 assign n_13 = ~n_22;
 assign n_21 = ~n_22;
 assign n_22 = ~n_20;
 assign n_20 = ~n_38;
 assign n_38 = ~in2_10_32_;
 assign in2_2 = ((in2_1_0_ & ~in2_1_32_) | ({in2[5]} & in2_1_32_));
 assign in2_5_1_ = ((in2_4_1_ & ~in2_4_32_) | (in2_2 & in2_4_32_));
 assign in2_5_0_ = ((in2_4_0_ & ~in2_4_32_) | ({in2[4]} & in2_4_32_));
 assign in2_8_2_ = ((in2_7_2_ & ~in2_7_32_) | (in2_5_1_ & in2_7_32_));
 assign in2_8_1_ = ((in2_7_1_ & ~in2_7_32_) | (in2_5_0_ & in2_7_32_));
 assign in2_8_0_ = ((in2_7_0_ & ~in2_7_32_) | ({in2[3]} & in2_7_32_));
 assign {out1[5]} = ((in2_16_5_ & ~in2_16_32_) | (in2_14_4_ & in2_16_32_));
 assign {out1[2]} = ((in2_16_2_ & ~in2_16_32_) | (in2_14_1_ & in2_16_32_));
 assign {out1[1]} = ((in2_16_1_ & ~in2_16_32_) | (in2_14_0_ & in2_16_32_));
 assign {out1[4]} = ((in2_16_4_ & ~in2_16_32_) | (in2_14_3_ & in2_16_32_));
 assign {out1[3]} = ((in2_16_3_ & ~in2_16_32_) | (in2_14_2_ & in2_16_32_));
 assign in2_10_32_ = ~(((sub_115_2_n_25 & sub_115_2_n_20) & ~{in1[10]}) & ~{in1[11]});
 assign sub_115_2_n_25 = ~(({in1[8]} | {in1[9]}) | sub_115_2_n_24);
 assign sub_115_2_n_24 = ~(((sub_115_2_n_23 & sub_115_2_n_10) & ~{in1[5]}) & ~{in1[6]});
 assign sub_115_2_n_23 = ~(({in1[7]} | {in1[4]}) | (sub_115_2_n_21 & sub_115_2_n_3));
 assign in2_10_3_ = ~(sub_115_2_n_13 ^ sub_115_2_n_19);
 assign sub_115_2_n_21 = ~(sub_115_2_n_2 & (sub_115_2_n_7 | (sub_115_2_n_16 & sub_115_2_n_6)));
 assign sub_115_2_n_20 = ~(({in1[22]} | {in1[23]}) | sub_115_2_n_17);
 assign sub_115_2_n_19 = (sub_115_2_n_7 | (sub_115_2_n_16 & sub_115_2_n_6));
 assign in2_10_2_ = ~(sub_115_2_n_12 ^ sub_115_2_n_16);
 assign sub_115_2_n_17 = ~(((sub_115_2_n_14 & sub_115_2_n_8) & ~{in1[20]}) & ~{in1[21]});
 assign sub_115_2_n_16 = ((sub_115_2_n_1 & sub_115_2_n_4) | (in2_8_0_ & (sub_115_2_n_1 ^ sub_115_2_n_4)));
 assign in2_10_1_ = ((in2_8_0_ ^ sub_115_2_n_1) ^ sub_115_2_n_4);
 assign sub_115_2_n_14 = ~((({in1[30]} | {in1[29]}) | ~sub_115_2_n_9) | ~sub_115_2_n_5);
 assign sub_115_2_n_13 = ~(sub_115_2_n_3 & sub_115_2_n_2);
 assign sub_115_2_n_12 = ~(~sub_115_2_n_7 & sub_115_2_n_6);
 assign in2_10_0_ = ~(sub_115_2_n_4 & (~{in2[2]} | {in1[0]}));
 assign sub_115_2_n_10 = ~((({in1[12]} | {in1[13]}) | {in1[14]}) | {in1[15]});
 assign sub_115_2_n_9 = ~((({in1[24]} | {in1[25]}) | {in1[26]}) | {in1[27]});
 assign sub_115_2_n_8 = ~((({in1[16]} | {in1[17]}) | {in1[18]}) | {in1[19]});
 assign sub_115_2_n_7 = ~(~in2_8_1_ | {in1[2]});
 assign sub_115_2_n_6 = ~(~in2_8_1_ & {in1[2]});
 assign sub_115_2_n_5 = ~({in1[28]} | {in1[31]});
 assign sub_115_2_n_4 = ~(~{in2[2]} & {in1[0]});
 assign sub_115_2_n_3 = ~(~{in1[3]} & in2_8_2_);
 assign sub_115_2_n_2 = ~(~in2_8_2_ & {in1[3]});
 assign sub_115_2_n_1 = ~{in1[1]};
 assign sub_134_2_n_31 = ~(sub_134_2_n_29 & ((sub_134_2_n_2 | sub_134_2_n_3) | {in1[5]}));
 assign sub_134_2_n_29 = (((sub_134_2_n_28 | sub_134_2_n_2) | sub_134_2_n_12) | {in1[5]});
 assign sub_134_2_n_28 = ~(sub_134_2_n_11 | (sub_134_2_n_0 & sub_134_2_n_10));
 assign sub_134_2_n_24 = ~(((sub_134_2_n_23 & sub_134_2_n_14) & ~{in1[16]}) & ~{in1[17]});
 assign sub_134_2_n_23 = ~((({in1[30]} | {in1[29]}) | ~sub_134_2_n_13) | ~sub_134_2_n_8);
 assign sub_134_2_n_22 = ~(sub_134_2_n_6 | (sub_134_2_n_4 & sub_134_2_n_5));
 assign sub_134_2_n_20 = ~(sub_134_2_n_12 | ~sub_134_2_n_3);
 assign sub_134_2_n_19 = ~(~sub_134_2_n_11 & sub_134_2_n_10);
 assign sub_134_2_n_18 = ~(sub_134_2_n_7 | ~sub_134_2_n_9);
 assign sub_134_2_n_17 = ~(~sub_134_2_n_6 & sub_134_2_n_5);
 assign sub_134_2_n_15 = ~((({in1[8]} | {in1[9]}) | {in1[10]}) | {in1[11]});
 assign sub_134_2_n_14 = ~((({in1[20]} | {in1[21]}) | {in1[22]}) | {in1[23]});
 assign sub_134_2_n_13 = ~((({in1[24]} | {in1[25]}) | {in1[26]}) | {in1[27]});
 assign sub_134_2_n_12 = ~(~{in1[4]} | in2_11_3_);
 assign sub_134_2_n_11 = ~({in1[3]} | ~in2_11_2_);
 assign sub_134_2_n_10 = ~(~in2_11_2_ & {in1[3]});
 assign sub_134_2_n_9 = ~(~{in1[2]} & in2_11_1_);
 assign sub_134_2_n_8 = ~({in1[28]} | {in1[31]});
 assign sub_134_2_n_7 = ~(~{in1[2]} | in2_11_1_);
 assign sub_134_2_n_6 = ~({in1[1]} | ~in2_11_0_);
 assign sub_134_2_n_5 = ~(~in2_11_0_ & {in1[1]});
 assign sub_134_2_n_4 = ~(~{in2[1]} & {in1[0]});
 assign sub_134_2_n_3 = ~(~{in1[4]} & in2_11_3_);
 assign sub_134_2_n_2 = ({in1[6]} | {in1[7]});
 assign sub_134_2_n_0 = ~(sub_134_2_n_9 & (sub_134_2_n_22 | sub_134_2_n_7));
 assign in2_16_5_ = ~(sub_153_2_n_22 ^ sub_153_2_n_35);
 assign sub_153_2_n_35 = ~(sub_153_2_n_2 & (sub_153_2_n_32 | sub_153_2_n_14));
 assign in2_16_4_ = ~(sub_153_2_n_20 ^ sub_153_2_n_32);
 assign sub_153_2_n_32 = ~(sub_153_2_n_13 | (sub_153_2_n_0 & sub_153_2_n_11));
 assign in2_16_3_ = ~(sub_153_2_n_19 ^ sub_153_2_n_0);
 assign in2_16_2_ = ~(sub_153_2_n_26 ^ sub_153_2_n_23);
 assign sub_153_2_n_28 = ~(((sub_153_2_n_27 & sub_153_2_n_16) & ~{in1[20]}) & ~{in1[21]});
 assign sub_153_2_n_27 = ~((({in1[30]} | {in1[29]}) | ~sub_153_2_n_15) | ~sub_153_2_n_12);
 assign sub_153_2_n_24 = ~(sub_153_2_n_5 & (~sub_153_2_n_3 | sub_153_2_n_2));
 assign sub_153_2_n_23 = ~(sub_153_2_n_9 | ~sub_153_2_n_10);
 assign sub_153_2_n_22 = ~(sub_153_2_n_5 & sub_153_2_n_3);
 assign sub_153_2_n_21 = ~(~sub_153_2_n_8 & sub_153_2_n_7);
 assign sub_153_2_n_20 = ~(sub_153_2_n_14 | ~sub_153_2_n_2);
 assign sub_153_2_n_19 = ~(~sub_153_2_n_13 & sub_153_2_n_11);
 assign sub_153_2_n_16 = ~((({in1[16]} | {in1[17]}) | {in1[18]}) | {in1[19]});
 assign sub_153_2_n_15 = ~((({in1[24]} | {in1[25]}) | {in1[26]}) | {in1[27]});
 assign sub_153_2_n_12 = ~({in1[28]} | {in1[31]});
 assign sub_153_2_n_0 = ~(sub_153_2_n_10 & (sub_153_2_n_26 | sub_153_2_n_9));
 assign in2_1_32_ = ~(((sub_58_2_n_12 & sub_58_2_n_11) & ~{in1[8]}) & ~{in1[9]});
 assign sub_58_2_n_12 = ~((({in1[10]} | {in1[11]}) | ~sub_58_2_n_10) | ~sub_58_2_n_5);
 assign sub_58_2_n_11 = ~(({in1[26]} | {in1[27]}) | sub_58_2_n_9);
 assign sub_58_2_n_10 = ~(((~sub_58_2_n_8 | {in1[7]}) | {in1[5]}) | {in1[6]});
 assign sub_58_2_n_9 = ~(((sub_58_2_n_7 & sub_58_2_n_4) & ~{in1[24]}) & ~{in1[25]});
 assign sub_58_2_n_8 = ~(((~sub_58_2_n_6 | {in1[2]}) | {in1[3]}) | {in1[4]});
 assign sub_58_2_n_7 = ~((({in1[20]} | {in1[23]}) | ~sub_58_2_n_3) | ~sub_58_2_n_1);
 assign sub_58_2_n_6 = ~({in1[1]} | (~{in2[5]} & {in1[0]}));
 assign sub_58_2_n_5 = ~((({in1[12]} | {in1[13]}) | {in1[14]}) | {in1[15]});
 assign sub_58_2_n_4 = ~((({in1[28]} | {in1[29]}) | {in1[30]}) | {in1[31]});
 assign sub_58_2_n_3 = ~((({in1[16]} | {in1[17]}) | {in1[18]}) | {in1[19]});
 assign in2_1_0_ = ({in1[0]} ^ {in2[5]});
 assign sub_58_2_n_1 = ~({in1[21]} | {in1[22]});
 assign in2_4_32_ = ~(((sub_77_2_n_17 & sub_77_2_n_14) & ~{in1[10]}) & ~{in1[11]});
 assign sub_77_2_n_17 = ~((({in1[8]} | {in1[9]}) | ~sub_77_2_n_16) | ~sub_77_2_n_7);
 assign sub_77_2_n_16 = ~(((~sub_77_2_n_15 | {in1[5]}) | {in1[4]}) | {in1[7]});
 assign sub_77_2_n_15 = ~((({in1[2]} | {in1[3]}) | sub_77_2_n_11) | {in1[6]});
 assign sub_77_2_n_14 = ~(({in1[26]} | {in1[27]}) | sub_77_2_n_13);
 assign sub_77_2_n_13 = ~(((sub_77_2_n_12 & sub_77_2_n_6) & ~{in1[24]}) & ~{in1[25]});
 assign sub_77_2_n_12 = ~((({in1[16]} | {in1[19]}) | ~sub_77_2_n_5) | ~sub_77_2_n_2);
 assign sub_77_2_n_11 = ~(sub_77_2_n_1 | (sub_77_2_n_4 & sub_77_2_n_3));
 assign in2_4_1_ = ~(sub_77_2_n_4 ^ sub_77_2_n_9);
 assign sub_77_2_n_9 = ~(~sub_77_2_n_1 & sub_77_2_n_3);
 assign in2_4_0_ = ~(sub_77_2_n_4 & (~{in2[4]} | {in1[0]}));
 assign sub_77_2_n_7 = ~((({in1[12]} | {in1[13]}) | {in1[14]}) | {in1[15]});
 assign sub_77_2_n_6 = ~((({in1[28]} | {in1[29]}) | {in1[30]}) | {in1[31]});
 assign sub_77_2_n_5 = ~((({in1[20]} | {in1[21]}) | {in1[22]}) | {in1[23]});
 assign sub_77_2_n_4 = ~(~{in2[4]} & {in1[0]});
 assign sub_77_2_n_3 = ~(~in2_2 & {in1[1]});
 assign sub_77_2_n_2 = ~({in1[17]} | {in1[18]});
 assign sub_77_2_n_1 = ~({in1[1]} | ~in2_2);
 assign in2_7_32_ = ~(((sub_96_2_n_20 & sub_96_2_n_17) & ~{in1[10]}) & ~{in1[11]});
 assign sub_96_2_n_20 = ~(({in1[8]} | {in1[9]}) | sub_96_2_n_19);
 assign sub_96_2_n_19 = ~(((sub_96_2_n_18 & sub_96_2_n_8) & ~{in1[5]}) & ~{in1[6]});
 assign sub_96_2_n_18 = ~(((sub_96_2_n_16 | {in1[3]}) | {in1[4]}) | {in1[7]});
 assign sub_96_2_n_17 = ~(({in1[18]} | {in1[19]}) | sub_96_2_n_14);
 assign sub_96_2_n_16 = ~(sub_96_2_n_2 | (sub_96_2_n_13 & sub_96_2_n_5));
 assign in2_7_2_ = ~(sub_96_2_n_10 ^ sub_96_2_n_13);
 assign sub_96_2_n_14 = ~(((sub_96_2_n_11 & sub_96_2_n_7) & ~{in1[16]}) & ~{in1[17]});
 assign sub_96_2_n_13 = ((sub_96_2_n_1 & sub_96_2_n_3) | (in2_5_0_ & (sub_96_2_n_1 ^ sub_96_2_n_3)));
 assign in2_7_1_ = ((in2_5_0_ ^ sub_96_2_n_1) ^ sub_96_2_n_3);
 assign sub_96_2_n_11 = ~((({in1[26]} | {in1[25]}) | ~sub_96_2_n_6) | ~sub_96_2_n_4);
 assign sub_96_2_n_10 = ~(~sub_96_2_n_2 & sub_96_2_n_5);
 assign in2_7_0_ = ~(sub_96_2_n_3 & (~{in2[3]} | {in1[0]}));
 assign sub_96_2_n_8 = ~((({in1[12]} | {in1[13]}) | {in1[14]}) | {in1[15]});
 assign sub_96_2_n_7 = ~((({in1[20]} | {in1[21]}) | {in1[22]}) | {in1[23]});
 assign sub_96_2_n_6 = ~((({in1[28]} | {in1[29]}) | {in1[30]}) | {in1[31]});
 assign sub_96_2_n_5 = ~(~in2_5_1_ & {in1[2]});
 assign sub_96_2_n_4 = ~({in1[24]} | {in1[27]});
 assign sub_96_2_n_3 = ~(~{in2[3]} & {in1[0]});
 assign sub_96_2_n_2 = ~({in1[2]} | ~in2_5_1_);
 assign sub_96_2_n_1 = ~{in1[1]};
 assign n_104 = ~((n_34 & ~stall) | (n_80 & stall));
assign out1[6] = 1'B0;
endmodule
